module Gowin_MIPI_DPHY_RX (d0ln_hsrxd, d1ln_hsrxd, d0ln_hsrxd_vld, d1ln_hsrxd_vld, di_lprx0_n, di_lprx0_p, di_lprx1_n, di_lprx1_p, di_lprxck_n, di_lprxck_p, rx_clk_o, deskew_error, d0ln_deskew_done, d1ln_deskew_done, ck_n, ck_p, rx0_n, rx0_p, rx1_n, rx1_p, lprx_en_ck, lprx_en_d0, lprx_en_d1, hsrx_odten_ck, hsrx_odten_d0, hsrx_odten_d1, d0ln_hsrx_dren, d1ln_hsrx_dren, hsrx_en_ck, hs_8bit_mode, rx_clk_1x, rx_invert, lalign_en, walign_by, do_lptx0_n, do_lptx0_p, do_lptx1_n, do_lptx1_p, do_lptxck_n, do_lptxck_p, lptx_en_ck, lptx_en_d0, lptx_en_d1, byte_lendian, hsrx_stop, pwron, reset, deskew_lnsel, deskew_mth, deskew_owval, deskew_req, drst_n, one_byte0_match, word_lendian, fifo_rd_std, deskew_by, deskew_en_oedge, deskew_half_opening, deskew_lsb_mode, deskew_m, deskew_mset, deskew_oclkedg_en, eqcs_lane0, eqcs_lane1, eqcs_ck, eqrs_lane0, eqrs_lane1, eqrs_ck, hsrx_dlydir_lane0, hsrx_dlydir_lane1, hsrx_dlydir_ck, hsrx_dlyldn_lane0, hsrx_dlyldn_lane1, hsrx_dlyldn_ck, hsrx_dlymv_lane0, hsrx_dlymv_lane1, hsrx_dlymv_ck, walign_dvld);

output [15:0] d0ln_hsrxd;
output [15:0] d1ln_hsrxd;
output d0ln_hsrxd_vld;
output d1ln_hsrxd_vld;
output di_lprx0_n;
output di_lprx0_p;
output di_lprx1_n;
output di_lprx1_p;
output di_lprxck_n;
output di_lprxck_p;
output rx_clk_o;
output deskew_error;
output d0ln_deskew_done;
output d1ln_deskew_done;
inout ck_n;
inout ck_p;
inout rx0_n;
inout rx0_p;
inout rx1_n;
inout rx1_p;
input lprx_en_ck;
input lprx_en_d0;
input lprx_en_d1;
input hsrx_odten_ck;
input hsrx_odten_d0;
input hsrx_odten_d1;
input d0ln_hsrx_dren;
input d1ln_hsrx_dren;
input hsrx_en_ck;
input hs_8bit_mode;
input rx_clk_1x;
input rx_invert;
input lalign_en;
input walign_by;
input do_lptx0_n;
input do_lptx0_p;
input do_lptx1_n;
input do_lptx1_p;
input do_lptxck_n;
input do_lptxck_p;
input lptx_en_ck;
input lptx_en_d0;
input lptx_en_d1;
input byte_lendian;
input hsrx_stop;
input pwron;
input reset;
input [2:0] deskew_lnsel;
input [12:0] deskew_mth;
input [6:0] deskew_owval;
input deskew_req;
input drst_n;
input one_byte0_match;
input word_lendian;
input [2:0] fifo_rd_std;
input deskew_by;
input deskew_en_oedge;
input [5:0] deskew_half_opening;
input [1:0] deskew_lsb_mode;
input [2:0] deskew_m;
input [6:0] deskew_mset;
input deskew_oclkedg_en;
input [2:0] eqcs_lane0;
input [2:0] eqcs_lane1;
input [2:0] eqcs_ck;
input [2:0] eqrs_lane0;
input [2:0] eqrs_lane1;
input [2:0] eqrs_ck;
input hsrx_dlydir_lane0;
input hsrx_dlydir_lane1;
input hsrx_dlydir_ck;
input hsrx_dlyldn_lane0;
input hsrx_dlyldn_lane1;
input hsrx_dlyldn_ck;
input hsrx_dlymv_lane0;
input hsrx_dlymv_lane1;
input hsrx_dlymv_ck;
input walign_dvld;

wire [15:0] d2ln_hsrxd;
wire [15:0] d3ln_hsrxd;
wire d2ln_hsrxd_vld;
wire d3ln_hsrxd_vld;
wire di_lprx2_n;
wire di_lprx2_p;
wire di_lprx3_n;
wire di_lprx3_p;
wire d2ln_deskew_done;
wire d3ln_deskew_done;
wire rx2_n;
wire rx2_p;
wire rx3_n;
wire rx3_p;
wire gw_gnd;

endmodule

