


`timescale 1ns / 1ps
`default_nettype none


module top
		#(
			parameter	X_WIDTH   = 10,
			parameter	Y_WIDTH   = 8,
			parameter	X_NUM     = 512,
			parameter	Y_NUM     = 128,
			parameter	MAX_X_NUM = 512,
			parameter	MAX_Y_NUM = 128
		)
		(
			input	wire			in_clk125,
			
			input	wire	[3:0]	push_sw,
			input	wire	[3:0]	dip_sw,
			output	wire	[3:0]	led,
			output	wire	[7:0]	pmod_a,
			
			input	wire			cam_clk_hs_p,
			input	wire			cam_clk_hs_n,
			input	wire			cam_clk_lp_p,
			input	wire			cam_clk_lp_n,
			input	wire	[1:0]	cam_data_hs_p,
			input	wire	[1:0]	cam_data_hs_n,
			input	wire	[1:0]	cam_data_lp_p,
			input	wire	[1:0]	cam_data_lp_n,
			input	wire			cam_clk,
			output	wire			cam_gpio,
			inout	wire			cam_scl,
			inout	wire			cam_sda,
			
			output	wire			hdmi_tx_clk_p,
			output	wire			hdmi_tx_clk_n,
			output	wire	[2:0]	hdmi_tx_data_p,
			output	wire	[2:0]	hdmi_tx_data_n,
			
			inout	wire	[14:0]	DDR_addr,
			inout	wire	[2:0]	DDR_ba,
			inout	wire			DDR_cas_n,
			inout	wire			DDR_ck_n,
			inout	wire			DDR_ck_p,
			inout	wire			DDR_cke,
			inout	wire			DDR_cs_n,
			inout	wire	[3:0]	DDR_dm,
			inout	wire	[31:0]	DDR_dq,
			inout	wire	[3:0]	DDR_dqs_n,
			inout	wire	[3:0]	DDR_dqs_p,
			inout	wire			DDR_odt,
			inout	wire			DDR_ras_n,
			inout	wire			DDR_reset_n,
			inout	wire			DDR_we_n,
			inout	wire			FIXED_IO_ddr_vrn,
			inout	wire			FIXED_IO_ddr_vrp,
			inout	wire	[53:0]	FIXED_IO_mio,
			inout	wire			FIXED_IO_ps_clk,
			inout	wire			FIXED_IO_ps_porb,
			inout	wire			FIXED_IO_ps_srstb
		);
	
	
	// ----------------------------------------
	//  input clock
	// ----------------------------------------
	
	wire								in_clk125_i;
	wire								in_clk125_buf;
	IBUFG
		i_ibufg_in_clk125
			(
				.I	(in_clk125),
				.O	(in_clk125_i)
			);
	BUFG
		i_bufg_in_clk125
			(
				.I	(in_clk125_i),
				.O	(in_clk125_buf)
			);
	
	
	
	// ----------------------------------------
	//  block design (PS)
	// ----------------------------------------
	
						wire			sys_reset;
	(* KEEP = "true" *)	wire			sys_clk100;
	(* KEEP = "true" *)	wire			sys_clk200;
	(* KEEP = "true" *)	wire			sys_clk250;
	
						wire			vout_reset;
	(* KEEP = "true" *)	wire			vout_clk;
	(* KEEP = "true" *)	wire			vout_clk_x5;
	
	wire			axi4l_peri_aresetn;
	wire			axi4l_peri_aclk;
	wire	[31:0]	axi4l_peri_awaddr;
	wire	[2:0]	axi4l_peri_awprot;
	wire			axi4l_peri_awvalid;
	wire			axi4l_peri_awready;
	wire	[3:0]	axi4l_peri_wstrb;
	wire	[31:0]	axi4l_peri_wdata;
	wire			axi4l_peri_wvalid;
	wire			axi4l_peri_wready;
	wire	[1:0]	axi4l_peri_bresp;
	wire			axi4l_peri_bvalid;
	wire			axi4l_peri_bready;
	wire	[31:0]	axi4l_peri_araddr;
	wire	[2:0]	axi4l_peri_arprot;
	wire			axi4l_peri_arvalid;
	wire			axi4l_peri_arready;
	wire	[31:0]	axi4l_peri_rdata;
	wire	[1:0]	axi4l_peri_rresp;
	wire			axi4l_peri_rvalid;
	wire			axi4l_peri_rready;
	
	
	wire			axi4_mem_aresetn;
	wire			axi4_mem_aclk;
	
	wire	[5:0]	axi4_mem0_awid;
	wire	[31:0]	axi4_mem0_awaddr;
	wire	[1:0]	axi4_mem0_awburst;
	wire	[3:0]	axi4_mem0_awcache;
	wire	[7:0]	axi4_mem0_awlen;
	wire	[0:0]	axi4_mem0_awlock;
	wire	[2:0]	axi4_mem0_awprot;
	wire	[3:0]	axi4_mem0_awqos;
	wire	[3:0]	axi4_mem0_awregion;
	wire	[2:0]	axi4_mem0_awsize;
	wire			axi4_mem0_awvalid;
	wire			axi4_mem0_awready;
	wire	[7:0]	axi4_mem0_wstrb;
	wire	[63:0]	axi4_mem0_wdata;
	wire			axi4_mem0_wlast;
	wire			axi4_mem0_wvalid;
	wire			axi4_mem0_wready;
	wire	[5:0]	axi4_mem0_bid;
	wire	[1:0]	axi4_mem0_bresp;
	wire			axi4_mem0_bvalid;
	wire			axi4_mem0_bready;
	wire	[5:0]	axi4_mem0_arid;
	wire	[31:0]	axi4_mem0_araddr;
	wire	[1:0]	axi4_mem0_arburst;
	wire	[3:0]	axi4_mem0_arcache;
	wire	[7:0]	axi4_mem0_arlen;
	wire	[0:0]	axi4_mem0_arlock;
	wire	[2:0]	axi4_mem0_arprot;
	wire	[3:0]	axi4_mem0_arqos;
	wire	[3:0]	axi4_mem0_arregion;
	wire	[2:0]	axi4_mem0_arsize;
	wire			axi4_mem0_arvalid;
	wire			axi4_mem0_arready;
	wire	[5:0]	axi4_mem0_rid;
	wire	[1:0]	axi4_mem0_rresp;
	wire	[63:0]	axi4_mem0_rdata;
	wire			axi4_mem0_rlast;
	wire			axi4_mem0_rvalid;
	wire			axi4_mem0_rready;
	
	wire			IIC_0_0_scl_i;
	wire			IIC_0_0_scl_o;
	wire			IIC_0_0_scl_t;
	wire			IIC_0_0_sda_i;
	wire			IIC_0_0_sda_o;
	wire			IIC_0_0_sda_t;
	
	design_1
		i_design_1
			(
				.sys_reset				(1'b0),
				.sys_clock				(in_clk125_buf),
				
				.out_reset				(sys_reset),
				.out_clk100				(sys_clk100),
				.out_clk200				(sys_clk200),
				.out_clk250				(sys_clk250),
				
				.vout_reset				(vout_reset),
				.vout_clk				(vout_clk),
				.vout_clk_x5			(vout_clk_x5),
				
				.m_axi4l_peri_aresetn	(axi4l_peri_aresetn),
				.m_axi4l_peri_aclk		(axi4l_peri_aclk),
				.m_axi4l_peri_awaddr	(axi4l_peri_awaddr),
				.m_axi4l_peri_awprot	(axi4l_peri_awprot),
				.m_axi4l_peri_awvalid	(axi4l_peri_awvalid),
				.m_axi4l_peri_awready	(axi4l_peri_awready),
				.m_axi4l_peri_wstrb		(axi4l_peri_wstrb),
				.m_axi4l_peri_wdata		(axi4l_peri_wdata),
				.m_axi4l_peri_wvalid	(axi4l_peri_wvalid),
				.m_axi4l_peri_wready	(axi4l_peri_wready),
				.m_axi4l_peri_bresp		(axi4l_peri_bresp),
				.m_axi4l_peri_bvalid	(axi4l_peri_bvalid),
				.m_axi4l_peri_bready	(axi4l_peri_bready),
				.m_axi4l_peri_araddr	(axi4l_peri_araddr),
				.m_axi4l_peri_arprot	(axi4l_peri_arprot),
				.m_axi4l_peri_arvalid	(axi4l_peri_arvalid),
				.m_axi4l_peri_arready	(axi4l_peri_arready),
				.m_axi4l_peri_rdata		(axi4l_peri_rdata),
				.m_axi4l_peri_rresp		(axi4l_peri_rresp),
				.m_axi4l_peri_rvalid	(axi4l_peri_rvalid),
				.m_axi4l_peri_rready	(axi4l_peri_rready),
				
				
				.s_axi4_mem_aresetn		(axi4_mem_aresetn),
				.s_axi4_mem_aclk		(axi4_mem_aclk),
				
				.s_axi4_mem0_awid		(axi4_mem0_awid),
				.s_axi4_mem0_awaddr		(axi4_mem0_awaddr),
				.s_axi4_mem0_awburst	(axi4_mem0_awburst),
				.s_axi4_mem0_awcache	(axi4_mem0_awcache),
				.s_axi4_mem0_awlen		(axi4_mem0_awlen),
				.s_axi4_mem0_awlock		(axi4_mem0_awlock),
				.s_axi4_mem0_awprot		(axi4_mem0_awprot),
				.s_axi4_mem0_awqos		(axi4_mem0_awqos),
	//			.s_axi4_mem0_awregion	(axi4_mem0_awregion),
				.s_axi4_mem0_awsize		(axi4_mem0_awsize),
				.s_axi4_mem0_awvalid	(axi4_mem0_awvalid),
				.s_axi4_mem0_awready	(axi4_mem0_awready),
				.s_axi4_mem0_wstrb		(axi4_mem0_wstrb),
				.s_axi4_mem0_wdata		(axi4_mem0_wdata),
				.s_axi4_mem0_wlast		(axi4_mem0_wlast),
				.s_axi4_mem0_wvalid		(axi4_mem0_wvalid),
				.s_axi4_mem0_wready		(axi4_mem0_wready),
				.s_axi4_mem0_bid		(axi4_mem0_bid),
				.s_axi4_mem0_bresp		(axi4_mem0_bresp),
				.s_axi4_mem0_bvalid		(axi4_mem0_bvalid),
				.s_axi4_mem0_bready		(axi4_mem0_bready),
				.s_axi4_mem0_araddr		(axi4_mem0_araddr),
				.s_axi4_mem0_arburst	(axi4_mem0_arburst),
				.s_axi4_mem0_arcache	(axi4_mem0_arcache),
				.s_axi4_mem0_arid		(axi4_mem0_arid),
				.s_axi4_mem0_arlen		(axi4_mem0_arlen),
				.s_axi4_mem0_arlock		(axi4_mem0_arlock),
				.s_axi4_mem0_arprot		(axi4_mem0_arprot),
				.s_axi4_mem0_arqos		(axi4_mem0_arqos),
	//			.s_axi4_mem0_arregion	(axi4_mem0_arregion),
				.s_axi4_mem0_arsize		(axi4_mem0_arsize),
				.s_axi4_mem0_arvalid	(axi4_mem0_arvalid),
				.s_axi4_mem0_arready	(axi4_mem0_arready),
				.s_axi4_mem0_rid		(axi4_mem0_rid),
				.s_axi4_mem0_rresp		(axi4_mem0_rresp),
				.s_axi4_mem0_rdata		(axi4_mem0_rdata),
				.s_axi4_mem0_rlast		(axi4_mem0_rlast),
				.s_axi4_mem0_rvalid		(axi4_mem0_rvalid),
				.s_axi4_mem0_rready		(axi4_mem0_rready),
				
				.DDR_addr				(DDR_addr),
				.DDR_ba					(DDR_ba),
				.DDR_cas_n				(DDR_cas_n),
				.DDR_ck_n				(DDR_ck_n),
				.DDR_ck_p				(DDR_ck_p),
				.DDR_cke				(DDR_cke),
				.DDR_cs_n				(DDR_cs_n),
				.DDR_dm					(DDR_dm),
				.DDR_dq					(DDR_dq),
				.DDR_dqs_n				(DDR_dqs_n),
				.DDR_dqs_p				(DDR_dqs_p),
				.DDR_odt				(DDR_odt),
				.DDR_ras_n				(DDR_ras_n),
				.DDR_reset_n			(DDR_reset_n),
				.DDR_we_n				(DDR_we_n),
				.FIXED_IO_ddr_vrn		(FIXED_IO_ddr_vrn),
				.FIXED_IO_ddr_vrp		(FIXED_IO_ddr_vrp),
				.FIXED_IO_mio			(FIXED_IO_mio),
				.FIXED_IO_ps_clk		(FIXED_IO_ps_clk),
				.FIXED_IO_ps_porb		(FIXED_IO_ps_porb),
				.FIXED_IO_ps_srstb		(FIXED_IO_ps_srstb),
				
				.IIC_0_0_scl_i			(IIC_0_0_scl_i),
				.IIC_0_0_scl_o			(IIC_0_0_scl_o),
				.IIC_0_0_scl_t			(IIC_0_0_scl_t),
				.IIC_0_0_sda_i			(IIC_0_0_sda_i),
				.IIC_0_0_sda_o			(IIC_0_0_sda_o),
				.IIC_0_0_sda_t			(IIC_0_0_sda_t)
			);
	
	assign cam_gpio = dip_sw[0];
	
	IOBUF
		i_IOBUF_cam_scl
			(
				.IO		(cam_scl),
				.I		(IIC_0_0_scl_o),
				.O		(IIC_0_0_scl_i),
				.T		(IIC_0_0_scl_t)
			);

	IOBUF
		i_iobuf_cam_sda
			(
				.IO		(cam_sda),
				.I		(IIC_0_0_sda_o),
				.O		(IIC_0_0_sda_i),
				.T		(IIC_0_0_sda_t)
			);
	
	
	// AXI4L => WISHBONE
								wire					wb_rst_o;
								wire					wb_clk_o;
	(* MARK_DEBUG = "true" *)	wire	[29:0]			wb_host_adr_o;
	(* MARK_DEBUG = "true" *)	wire	[31:0]			wb_host_dat_o;
	(* MARK_DEBUG = "true" *)	wire	[31:0]			wb_host_dat_i;
	(* MARK_DEBUG = "true" *)	wire					wb_host_we_o;
	(* MARK_DEBUG = "true" *)	wire	[3:0]			wb_host_sel_o;
	(* MARK_DEBUG = "true" *)	wire					wb_host_stb_o;
	(* MARK_DEBUG = "true" *)	wire					wb_host_ack_i;
	
	jelly_axi4l_to_wishbone
			#(
				.AXI4L_ADDR_WIDTH	(32),
				.AXI4L_DATA_SIZE	(2)		// 0:8bit, 1:16bit, 2:32bit ...
			)
		i_axi4l_to_wishbone
			(
				.s_axi4l_aresetn	(axi4l_peri_aresetn),
				.s_axi4l_aclk		(axi4l_peri_aclk),
				.s_axi4l_awaddr		(axi4l_peri_awaddr),
				.s_axi4l_awprot		(axi4l_peri_awprot),
				.s_axi4l_awvalid	(axi4l_peri_awvalid),
				.s_axi4l_awready	(axi4l_peri_awready),
				.s_axi4l_wstrb		(axi4l_peri_wstrb),
				.s_axi4l_wdata		(axi4l_peri_wdata),
				.s_axi4l_wvalid		(axi4l_peri_wvalid),
				.s_axi4l_wready		(axi4l_peri_wready),
				.s_axi4l_bresp		(axi4l_peri_bresp),
				.s_axi4l_bvalid		(axi4l_peri_bvalid),
				.s_axi4l_bready		(axi4l_peri_bready),
				.s_axi4l_araddr		(axi4l_peri_araddr),
				.s_axi4l_arprot		(axi4l_peri_arprot),
				.s_axi4l_arvalid	(axi4l_peri_arvalid),
				.s_axi4l_arready	(axi4l_peri_arready),
				.s_axi4l_rdata		(axi4l_peri_rdata),
				.s_axi4l_rresp		(axi4l_peri_rresp),
				.s_axi4l_rvalid		(axi4l_peri_rvalid),
				.s_axi4l_rready		(axi4l_peri_rready),
				
				.m_wb_rst_o			(wb_rst_o),
				.m_wb_clk_o			(wb_clk_o),
				.m_wb_adr_o			(wb_host_adr_o),
				.m_wb_dat_o			(wb_host_dat_o),
				.m_wb_dat_i			(wb_host_dat_i),
				.m_wb_we_o			(wb_host_we_o),
				.m_wb_sel_o			(wb_host_sel_o),
				.m_wb_stb_o			(wb_host_stb_o),
				.m_wb_ack_i			(wb_host_ack_i)
			);
	
	
	// ----------------------------------------
	//  Global ID
	// ----------------------------------------
	
	wire	[31:0]			wb_gid_dat_o;
	wire					wb_gid_stb_i;
	wire					wb_gid_ack_o;
	
	assign wb_gid_dat_o = 32'h01234567;
	assign wb_gid_ack_o = wb_gid_stb_i;
	
	
	
	// ----------------------------------------
	//  MIPI D-PHY RX
	// ----------------------------------------
	
	(* KEEP = "true" *)
	wire				rxbyteclkhs;
	wire				system_rst_out;
	wire				init_done;
	
	wire				cl_rxclkactivehs;
	wire				cl_stopstate;
	wire				cl_enable         = 1;
	wire				cl_rxulpsclknot;
	wire				cl_ulpsactivenot;
	
	wire	[7:0]		dl0_rxdatahs;
	wire				dl0_rxvalidhs;
	wire				dl0_rxactivehs;
	wire				dl0_rxsynchs;
	
	wire				dl0_forcerxmode   = 0;
	wire				dl0_stopstate;
	wire				dl0_enable        = 1;
	wire				dl0_ulpsactivenot;
	
	wire				dl0_rxclkesc;
	wire				dl0_rxlpdtesc;
	wire				dl0_rxulpsesc;
	wire	[3:0]		dl0_rxtriggeresc;
	wire	[7:0]		dl0_rxdataesc;
	wire				dl0_rxvalidesc;
	
	wire				dl0_errsoths;
	wire				dl0_errsotsynchs;
	wire				dl0_erresc;
	wire				dl0_errsyncesc;
	wire				dl0_errcontrol;
	
	wire	[7:0]		dl1_rxdatahs;
	wire				dl1_rxvalidhs;
	wire				dl1_rxactivehs;
	wire				dl1_rxsynchs;
	
	wire				dl1_forcerxmode   = 0;
	wire				dl1_stopstate;
	wire				dl1_enable        = 1;
	wire				dl1_ulpsactivenot;
	
	wire				dl1_rxclkesc;
	wire				dl1_rxlpdtesc;
	wire				dl1_rxulpsesc;
	wire	[3:0]		dl1_rxtriggeresc;
	wire	[7:0]		dl1_rxdataesc;
	wire				dl1_rxvalidesc;
	
	wire				dl1_errsoths;
	wire				dl1_errsotsynchs;
	wire				dl1_erresc;
	wire				dl1_errsyncesc;
	wire				dl1_errcontrol;
	
	
	reg		[31:0]		dbg_dl0_count;
	reg		[31:0]		dbg_dl1_count;
	always @(posedge rxbyteclkhs) begin
		if (dl0_rxactivehs ) begin
			dbg_dl0_count <= dbg_dl0_count + 1;
		end
		if ( dl0_rxsynchs ) begin
			dbg_dl0_count <= 0;
		end
		
		if (dl1_rxactivehs ) begin
			dbg_dl1_count <= dbg_dl1_count + 1;
		end
		if ( dl1_rxsynchs ) begin
			dbg_dl1_count <= 0;
		end
	end
	
	
	mipi_dphy_cam
		i_mipi_dphy_cam
			(
				.core_clk			(sys_clk200),
				.core_rst			(sys_reset),
				.rxbyteclkhs		(rxbyteclkhs),
				.system_rst_out		(system_rst_out),
				.init_done			(init_done),
				
				.cl_rxclkactivehs	(cl_rxclkactivehs),
				.cl_stopstate		(cl_stopstate),
				.cl_enable			(cl_enable),
				.cl_rxulpsclknot	(cl_rxulpsclknot),
				.cl_ulpsactivenot	(cl_ulpsactivenot),
				
				.dl0_rxdatahs		(dl0_rxdatahs),
				.dl0_rxvalidhs		(dl0_rxvalidhs),
				.dl0_rxactivehs		(dl0_rxactivehs),
				.dl0_rxsynchs		(dl0_rxsynchs),
				
				.dl0_forcerxmode	(dl0_forcerxmode),
				.dl0_stopstate		(dl0_stopstate),
				.dl0_enable			(dl0_enable),
				.dl0_ulpsactivenot	(dl0_ulpsactivenot),
				
				.dl0_rxclkesc		(dl0_rxclkesc),
				.dl0_rxlpdtesc		(dl0_rxlpdtesc),
				.dl0_rxulpsesc		(dl0_rxulpsesc),
				.dl0_rxtriggeresc	(dl0_rxtriggeresc),
				.dl0_rxdataesc		(dl0_rxdataesc),
				.dl0_rxvalidesc		(dl0_rxvalidesc),
				
				.dl0_errsoths		(dl0_errsoths),
				.dl0_errsotsynchs	(dl0_errsotsynchs),
				.dl0_erresc			(dl0_erresc),
				.dl0_errsyncesc		(dl0_errsyncesc),
				.dl0_errcontrol		(dl0_errcontrol),
				
				.dl1_rxdatahs		(dl1_rxdatahs),
				.dl1_rxvalidhs		(dl1_rxvalidhs),
				.dl1_rxactivehs		(dl1_rxactivehs),
				.dl1_rxsynchs		(dl1_rxsynchs),
				
				.dl1_forcerxmode	(dl1_forcerxmode),
				.dl1_stopstate		(dl1_stopstate),
				.dl1_enable			(dl1_enable),
				.dl1_ulpsactivenot	(dl1_ulpsactivenot),
				
				.dl1_rxclkesc		(dl1_rxclkesc),
				.dl1_rxlpdtesc		(dl1_rxlpdtesc),
				.dl1_rxulpsesc		(dl1_rxulpsesc),
				.dl1_rxtriggeresc	(dl1_rxtriggeresc),
				.dl1_rxdataesc		(dl1_rxdataesc),
				.dl1_rxvalidesc		(dl1_rxvalidesc),
				
				.dl1_errsoths		(dl1_errsoths),
				.dl1_errsotsynchs	(dl1_errsotsynchs),
				.dl1_erresc			(dl1_erresc),
				.dl1_errsyncesc		(dl1_errsyncesc),
				.dl1_errcontrol		(dl1_errcontrol),
				
				.clk_hs_rxp			(cam_clk_hs_p),
				.clk_hs_rxn			(cam_clk_hs_n),
				.clk_lp_rxp			(cam_clk_lp_p),
				.clk_lp_rxn			(cam_clk_lp_n),
				.data_hs_rxp		(cam_data_hs_p),
				.data_hs_rxn		(cam_data_hs_n),
				.data_lp_rxp		(cam_data_lp_p),
				.data_lp_rxn		(cam_data_lp_n)
		   );
	
	
//	wire		dphy_clk   = rxbyteclkhs;
//	wire		dphy_reset = system_rst_out;
	
	
	wire		dphy_clk   = rxbyteclkhs;
	wire		dphy_reset;
	jelly_reset
			#(
				.IN_LOW_ACTIVE		(0),
				.OUT_LOW_ACTIVE		(0),
				.INPUT_REGS			(2),
				.COUNTER_WIDTH		(5),
				.INSERT_BUFG		(0)
			)
		i_reset
			(
				.clk				(dphy_clk),
				.in_reset			(sys_reset || system_rst_out),
				.out_reset			(dphy_reset)
			);
	
	
	
	// ----------------------------------------
	//  CSI-2
	// ----------------------------------------
	
	wire			axi4s_cam_aresetn = ~sys_reset;
	wire			axi4s_cam_aclk    = sys_clk200;
	
	(* MARK_DEBUG = "true" *)	wire	[0:0]	axi4s_csi2_tuser;
	(* MARK_DEBUG = "true" *)	wire			axi4s_csi2_tlast;
	(* MARK_DEBUG = "true" *)	wire	[9:0]	axi4s_csi2_tdata;
	(* MARK_DEBUG = "true" *)	wire			axi4s_csi2_tvalid;
	(* MARK_DEBUG = "true" *)	wire			axi4s_csi2_tready;
	
	jelly_csi2_rx
			#(
				.LANE_NUM			(2),
				.DATA_WIDTH			(10),
				.M_FIFO_ASYNC		(1)
			)
		i_csi2_rx
			(
				.aresetn			(~sys_reset),
				.aclk				(sys_clk250),
				
				.rxreseths			(system_rst_out),
				.rxbyteclkhs		(rxbyteclkhs),
				.rxdatahs			({dl1_rxdatahs,   dl0_rxdatahs  }),
				.rxvalidhs			({dl1_rxvalidhs,  dl0_rxvalidhs }),
				.rxactivehs			({dl1_rxactivehs, dl0_rxactivehs}),
				.rxsynchs			({dl1_rxsynchs,   dl0_rxsynchs  }),
				
				.m_axi4s_aresetn	(axi4s_cam_aresetn),
				.m_axi4s_aclk		(axi4s_cam_aclk),
				.m_axi4s_tuser		(axi4s_csi2_tuser),
				.m_axi4s_tlast		(axi4s_csi2_tlast),
				.m_axi4s_tdata		(axi4s_csi2_tdata),
				.m_axi4s_tvalid		(axi4s_csi2_tvalid),
				.m_axi4s_tready		(1'b1)	// (axi4s_csi2_tready)
			);
	
	
	wire	[0:0]	axi4s_fifo_tuser;
	wire			axi4s_fifo_tlast;
	wire	[9:0]	axi4s_fifo_tdata;
	wire			axi4s_fifo_tvalid;
	wire			axi4s_fifo_tready;
	
	jelly_fifo_fwtf
			#(
				.DATA_WIDTH			(2+10),
				.PTR_WIDTH			(0),	// bypass
				.DOUT_REGS			(0),
				.RAM_TYPE			("block"),
				.LOW_DEALY			(0),
				.SLAVE_REGS			(0),
				.MASTER_REGS		(1)
			)
		i_fifo_fifo_fwtf_csi2
			(
				.reset				(~axi4s_cam_aresetn),
				.clk				(axi4s_cam_aclk),
				
				.s_data				({axi4s_csi2_tuser, axi4s_csi2_tlast, axi4s_csi2_tdata}),
				.s_valid			(axi4s_csi2_tvalid),
				.s_ready			(axi4s_csi2_tready),
				.s_free_count		(),
				
				.m_data				({axi4s_fifo_tuser, axi4s_fifo_tlast, axi4s_fifo_tdata}),
				.m_valid			(axi4s_fifo_tvalid),
				.m_ready			(axi4s_fifo_tready),
				.m_data_count		()
			);
	
	
	
	// normalize
	wire	[0:0]			axi4s_norm_tuser;
	wire					axi4s_norm_tlast;
	wire	[9:0]			axi4s_norm_tdata;
	wire					axi4s_norm_tvalid;
	wire					axi4s_norm_tready;
	
	wire	[31:0]			wb_norm_dat_o;
	wire					wb_norm_stb_i;
	wire					wb_norm_ack_o;
	
	wire	[X_WIDTH-1:0]	image_width;
	wire	[Y_WIDTH-1:0]	image_height;
	
	jelly_video_normalizer
			#(
				.WB_ADR_WIDTH		(8),
				.WB_DAT_WIDTH		(32),
				
				.TUSER_WIDTH		(1),
				.TDATA_WIDTH		(10),
				.X_WIDTH			(X_WIDTH),
				.Y_WIDTH			(Y_WIDTH),
				.TIMER_WIDTH		(32),
				.S_SLAVE_REGS		(1),
				.S_MASTER_REGS		(1),
				.M_SLAVE_REGS		(1),
				.M_MASTER_REGS		(1),
				
				.INIT_CONTROL		(2'b11),
				.INIT_SKIP			(1),
				.INIT_PARAM_WIDTH	(X_NUM),
				.INIT_PARAM_HEIGHT	(Y_NUM),
				.INIT_PARAM_FILL	(10'd0),
				.INIT_PARAM_TIMEOUT	(32'h00010000)
			)
		i_video_normalizer
			(
				.aresetn			(axi4s_cam_aresetn),
				.aclk				(axi4s_cam_aclk),
				.aclken				(1'b1),
				
				.s_wb_rst_i			(wb_rst_o),
				.s_wb_clk_i			(wb_clk_o),
				.s_wb_adr_i			(wb_host_adr_o[7:0]),
				.s_wb_dat_o			(wb_norm_dat_o),
				.s_wb_dat_i			(wb_host_dat_o),
				.s_wb_we_i			(wb_host_we_o),
				.s_wb_sel_i			(wb_host_sel_o),
				.s_wb_stb_i			(wb_norm_stb_i),
				.s_wb_ack_o			(wb_norm_ack_o),

				.out_param_width	(image_width),
				.out_param_height	(image_height),
				
				.s_axi4s_tuser		(axi4s_fifo_tuser),
				.s_axi4s_tlast		(axi4s_fifo_tlast),
				.s_axi4s_tdata		(axi4s_fifo_tdata),
				.s_axi4s_tvalid		(axi4s_fifo_tvalid),
				.s_axi4s_tready		(axi4s_fifo_tready),
				
				/*
				.s_axi4s_tuser		(axi4s_csi2_tuser),
				.s_axi4s_tlast		(axi4s_csi2_tlast),
				.s_axi4s_tdata		(axi4s_csi2_tdata),
				.s_axi4s_tvalid		(axi4s_csi2_tvalid),
				.s_axi4s_tready		(axi4s_csi2_tready),
				*/
				
				.m_axi4s_tuser		(axi4s_norm_tuser),
				.m_axi4s_tlast		(axi4s_norm_tlast),
				.m_axi4s_tdata		(axi4s_norm_tdata),
				.m_axi4s_tvalid		(axi4s_norm_tvalid),
				.m_axi4s_tready		(axi4s_norm_tready)
			);
	
	
	// ����
	wire	[0:0]		axi4s_rgb_tuser;
	wire				axi4s_rgb_tlast;
	wire	[39:0]		axi4s_rgb_tdata;
	wire				axi4s_rgb_tvalid;
	wire				axi4s_rgb_tready;
	
	wire	[31:0]		wb_rgb_dat_o;
	wire				wb_rgb_stb_i;
	wire				wb_rgb_ack_o;
	
	video_raw_to_rgb
			#(
				.WB_ADR_WIDTH		(10),
				.WB_DAT_WIDTH		(32),
				
				.DATA_WIDTH			(10),
				
				.IMG_Y_NUM			(Y_NUM),
				.IMG_Y_WIDTH		(Y_WIDTH),
				
				.TUSER_WIDTH		(1)
			)
		i_video_raw_to_rgb
			(
				.aresetn			(axi4s_cam_aresetn),
				.aclk				(axi4s_cam_aclk),
				
				.s_wb_rst_i			(wb_rst_o),
				.s_wb_clk_i			(wb_clk_o),
				.s_wb_adr_i			(wb_host_adr_o[9:0]),
				.s_wb_dat_o			(wb_rgb_dat_o),
				.s_wb_dat_i			(wb_host_dat_o),
				.s_wb_we_i			(wb_host_we_o),
				.s_wb_sel_i			(wb_host_sel_o),
				.s_wb_stb_i			(wb_rgb_stb_i),
				.s_wb_ack_o			(wb_rgb_ack_o),
				
				.s_axi4s_tuser		(axi4s_norm_tuser),
				.s_axi4s_tlast		(axi4s_norm_tlast),
				.s_axi4s_tdata		(axi4s_norm_tdata),
				.s_axi4s_tvalid		(axi4s_norm_tvalid),
				.s_axi4s_tready		(axi4s_norm_tready),
				
				.m_axi4s_tuser		(axi4s_rgb_tuser),
				.m_axi4s_tlast		(axi4s_rgb_tlast),
				.m_axi4s_tdata		(axi4s_rgb_tdata),
				.m_axi4s_tvalid		(axi4s_rgb_tvalid),
				.m_axi4s_tready		(axi4s_rgb_tready)
			);
	
	
	
	// ���m�N����
	wire	[23:0]		axi4s_rgb_trgb = {axi4s_rgb_tdata[29:22], axi4s_rgb_tdata[19:12], axi4s_rgb_tdata[9:2]};
	wire	[7:0]		axi4s_rgb_traw = axi4s_rgb_tdata[39:32];
	
	wire	[0:0]		axi4s_gray_tuser;
	wire				axi4s_gray_tlast;
	wire	[9:0]		axi4s_gray_tdata;
	wire				axi4s_gray_tvalid;
	
	jelly_video_rgb_to_gray
			#(
				.COMPONENT_NUM		(3),
				.DATA_WIDTH			(10),
				.TUSER_WIDTH		(1)
			)
		i_video_rgb_to_gray
			(
				.aresetn			(axi4s_cam_aresetn),
				.aclk				(axi4s_cam_aclk),
				
				.s_axi4s_tuser		(axi4s_rgb_tuser),
				.s_axi4s_tlast		(axi4s_rgb_tlast),
				.s_axi4s_tdata		(axi4s_rgb_tdata[29:0]),
				.s_axi4s_tvalid		(axi4s_rgb_tvalid),
				.s_axi4s_tready		(),
				
				.m_axi4s_tuser		(axi4s_gray_tuser),
				.m_axi4s_tlast		(axi4s_gray_tlast),
				.m_axi4s_tdata		(),
				.m_axi4s_tgray		(axi4s_gray_tdata),
				.m_axi4s_tvalid		(axi4s_gray_tvalid),
				.m_axi4s_tready		(1'b1)
			);
	
	
	// mnist
	wire	[0:0]			axi4s_mnist_tuser;
	wire					axi4s_mnist_tlast;
	wire	[3:0]			axi4s_mnist_tcount;
	wire	[3:0]			axi4s_mnist_tnumber;
	wire					axi4s_mnist_tvalid;
	
	wire	[31:0]			wb_mnist_dat_o;
	wire					wb_mnist_stb_i;
	wire					wb_mnist_ack_o;
	
	video_mnist
			#(
				.MAX_X_NUM			(MAX_X_NUM),
				.DATA_WIDTH			(8),
				.IMG_Y_NUM			(Y_NUM),
				.IMG_Y_WIDTH		(Y_WIDTH),
				.TUSER_WIDTH		(1),
				.WB_ADR_WIDTH		(10),
				.WB_DAT_WIDTH		(32),
				.INIT_PARAM_TH		(127),
				.INIT_PARAM_INV		(0)
			)
		i_video_mnist
			(
				.aresetn			(axi4s_cam_aresetn),
				.aclk				(axi4s_cam_aclk),
				
				.s_axi4s_tuser		(axi4s_gray_tuser),
				.s_axi4s_tlast		(axi4s_gray_tlast),
				.s_axi4s_tdata		(axi4s_gray_tdata[9:2]),
				.s_axi4s_tvalid		(axi4s_gray_tvalid),
				.s_axi4s_tready		(),
				
				.m_axi4s_tuser		(axi4s_mnist_tuser),
				.m_axi4s_tlast		(axi4s_mnist_tlast),
				.m_axi4s_tnumber	(axi4s_mnist_tnumber),
				.m_axi4s_tcount		(axi4s_mnist_tcount),
				.m_axi4s_tdata		(),
				.m_axi4s_tvalid		(axi4s_mnist_tvalid),
				.m_axi4s_tready		(1'b1),
				
				.s_wb_rst_i			(wb_rst_o),
				.s_wb_clk_i			(wb_clk_o),
				.s_wb_adr_i			(wb_host_adr_o[9:0]),
				.s_wb_dat_o			(wb_mnist_dat_o),
				.s_wb_dat_i			(wb_host_dat_o),
				.s_wb_we_i			(wb_host_we_o),
				.s_wb_sel_i			(wb_host_sel_o),
				.s_wb_stb_i			(wb_mnist_stb_i),
				.s_wb_ack_o			(wb_mnist_ack_o)
			);
	
	// frame buffer
	wire	[0:0]			axi4s_fmem_tuser;
	wire					axi4s_fmem_tlast;
	wire	[23:0]			axi4s_fmem_tdata;
	wire	[3:0]			axi4s_fmem_tcount;
	wire	[3:0]			axi4s_fmem_tnumber;
	wire					axi4s_fmem_tvalid;
	wire					axi4s_fmem_tready;
	
	video_dnn_fmem
			#(
				.TUSER_WIDTH			(1),
				.TDATA_WIDTH			(24),
				.STORE_TDATA_WIDTH		(4+4),
				
				.DIV_X					(2),
				.DIV_Y					(2),
				
				.X_WIDTH				(X_WIDTH),
				.Y_WIDTH				(Y_WIDTH),
				.MAX_X_NUM				(MAX_X_NUM),
				.MAX_Y_NUM				(MAX_Y_NUM),
				.RAM_TYPE				("block")
			)
		i_video_dnn_fmem
			(
				.aresetn				(axi4s_cam_aresetn),
				.aclk					(axi4s_cam_aclk),
				
				.s_axi4s_tuser			(axi4s_rgb_tuser),
				.s_axi4s_tlast			(axi4s_rgb_tlast),
				.s_axi4s_tdata			(axi4s_rgb_trgb),
				.s_axi4s_tvalid			(axi4s_rgb_tvalid),
				.s_axi4s_tready			(axi4s_rgb_tready),
				
				.m_axi4s_tuser			(axi4s_fmem_tuser),
				.m_axi4s_tlast			(axi4s_fmem_tlast),
				.m_axi4s_tdata			(axi4s_fmem_tdata),
				.m_axi4s_tdata_store	({axi4s_fmem_tnumber, axi4s_fmem_tcount}),
				.m_axi4s_tvalid			(axi4s_fmem_tvalid),
				.m_axi4s_tready			(axi4s_fmem_tready),
				
				
				.s_axi4s_store_aresetn	(axi4s_cam_aresetn),
				.s_axi4s_store_aclk		(axi4s_cam_aclk),
				.s_axi4s_store_tuser	(axi4s_mnist_tuser),
				.s_axi4s_store_tlast	(axi4s_mnist_tlast),
				.s_axi4s_store_tdata	({axi4s_mnist_tnumber, axi4s_mnist_tcount}),
				.s_axi4s_store_tvalid	(axi4s_mnist_tvalid)
			);
	
	
	// ���ʂŒ��F
	wire	[0:0]				axi4s_mcol_tuser;
	wire						axi4s_mcol_tlast;
	wire	[31:0]				axi4s_mcol_tdata;
	wire						axi4s_mcol_tvalid;
	wire						axi4s_mcol_tready;
	
	wire	[31:0]				wb_mcol_dat_o;
	wire						wb_mcol_stb_i;
	wire						wb_mcol_ack_o;
	
	video_mnist_color
			#(
				.DATA_WIDTH			(8),
				.TUSER_WIDTH		(1)
			)
		i_video_mnist_color
			(
				.aresetn			(axi4s_cam_aresetn),
				.aclk				(axi4s_cam_aclk),
				
				.s_axi4s_tuser		(axi4s_fmem_tuser),
				.s_axi4s_tlast		(axi4s_fmem_tlast),
				.s_axi4s_tnumber	(axi4s_fmem_tnumber),
				.s_axi4s_tcount		(axi4s_fmem_tcount),
				.s_axi4s_tdata		({8'h00, axi4s_fmem_tdata}),
				.s_axi4s_tbinary	(1'b0),
				.s_axi4s_tvalid		(axi4s_fmem_tvalid),
				.s_axi4s_tready		(axi4s_fmem_tready),
				
				.m_axi4s_tuser		(axi4s_mcol_tuser),
				.m_axi4s_tlast		(axi4s_mcol_tlast),
				.m_axi4s_tdata		(axi4s_mcol_tdata),
				.m_axi4s_tvalid		(axi4s_mcol_tvalid),
				.m_axi4s_tready		(axi4s_mcol_tready),
				
				.s_wb_rst_i			(wb_rst_o),
				.s_wb_clk_i			(wb_clk_o),
				.s_wb_adr_i			(wb_host_adr_o[7:0]),
				.s_wb_dat_o			(wb_mcol_dat_o),
				.s_wb_dat_i			(wb_host_dat_o),
				.s_wb_we_i			(wb_host_we_o),
				.s_wb_sel_i			(wb_host_sel_o),
				.s_wb_stb_i			(wb_mcol_stb_i),
				.s_wb_ack_o			(wb_mcol_ack_o)
			);
	
	
	
	// integrator
	wire	[0:0]				axi4s_int_tuser;
	wire						axi4s_int_tlast;
	wire	[23:0]				axi4s_int_tdata;
	wire						axi4s_int_tvalid;
	wire						axi4s_int_tready;
	
	wire	[31:0]				wb_int_dat_o;
	wire						wb_int_stb_i;
	wire						wb_int_ack_o;
	
	jelly_video_integrator_bram
			#(
				.COMPONENT_NUM			(3),
				.DATA_WIDTH				(8),
				.RATE_WIDTH				(8),
				.WB_ADR_WIDTH			(8),
				.WB_DAT_WIDTH			(32),
				.TUSER_WIDTH			(1),
				.X_WIDTH				(9),
				.Y_WIDTH				(8),
				.MAX_X_NUM				(512),
				.MAX_Y_NUM				(128),
				.RAM_TYPE				("block"),
				.FILLMEM				(1),
				.FILLMEM_DATA			(24'h7f7f7f),
				.COMPACT				(0),
				.ROUNDING				(1),
				.INIT_PARAM_RATE		(8'hf0)
			)
		i_video_integrator_bram
			(
				.aresetn				(axi4s_cam_aresetn),
				.aclk					(axi4s_cam_aclk),
				.aclken					(1'b1),
				
				.s_wb_rst_i				(wb_rst_o),
				.s_wb_clk_i				(wb_clk_o),
				.s_wb_adr_i				(wb_host_adr_o[7:0]),
				.s_wb_dat_o				(wb_int_dat_o),
				.s_wb_dat_i				(wb_host_dat_o),
				.s_wb_we_i				(wb_host_we_o),
				.s_wb_sel_i				(wb_host_sel_o),
				.s_wb_stb_i				(wb_int_stb_i),
				.s_wb_ack_o				(wb_int_ack_o),
				
				.s_axi4s_tuser			(axi4s_mcol_tuser),
				.s_axi4s_tlast			(axi4s_mcol_tlast),
				.s_axi4s_tdata			(axi4s_mcol_tdata[23:0]),
				.s_axi4s_tvalid			(axi4s_mcol_tvalid),
				.s_axi4s_tready			(axi4s_mcol_tready),
				
				.m_axi4s_tuser			(axi4s_int_tuser),
				.m_axi4s_tlast			(axi4s_int_tlast),
				.m_axi4s_tdata			(axi4s_int_tdata),
				.m_axi4s_tvalid			(axi4s_int_tvalid),
				.m_axi4s_tready			(axi4s_int_tready)
			);
	
	
	// DMA write
	wire	[31:0]			wb_vdmaw_dat_o;
	wire					wb_vdmaw_stb_i;
	wire					wb_vdmaw_ack_o;
	
	jelly_vdma_axi4s_to_axi4
			#(
				.ASYNC				(1),
				.FIFO_PTR_WIDTH		(12),
				
				.PIXEL_SIZE			(2),	// 32bit
				.AXI4_ID_WIDTH		(6),
				.AXI4_ADDR_WIDTH	(32),
				.AXI4_DATA_SIZE		(3),	// 64bit
				.AXI4S_DATA_SIZE	(2),	// 32bit
				.AXI4S_USER_WIDTH	(1),
				.INDEX_WIDTH		(8),
				.STRIDE_WIDTH		(16),
				.H_WIDTH			(14),
				.V_WIDTH			(14),
				.SIZE_WIDTH			(32),
				
				.WB_ADR_WIDTH		(8),
				.WB_DAT_WIDTH		(32),
				
				.INIT_CTL_CONTROL	(2'b00),
				.INIT_PARAM_ADDR	(32'h3000_0000),
//				.INIT_PARAM_STRIDE	(X_NUM*2),
				.INIT_PARAM_STRIDE	(8192),
				.INIT_PARAM_WIDTH	(X_NUM),
				.INIT_PARAM_HEIGHT	(Y_NUM),
				.INIT_PARAM_SIZE	(X_NUM*Y_NUM),
				.INIT_PARAM_AWLEN	(7)
			)
		i_vdma_axi4s_to_axi4
			(
				.m_axi4_aresetn		(axi4_mem_aresetn),
				.m_axi4_aclk		(axi4_mem_aclk),
				.m_axi4_awid		(axi4_mem0_awid),
				.m_axi4_awaddr		(axi4_mem0_awaddr),
				.m_axi4_awburst		(axi4_mem0_awburst),
				.m_axi4_awcache		(axi4_mem0_awcache),
				.m_axi4_awlen		(axi4_mem0_awlen),
				.m_axi4_awlock		(axi4_mem0_awlock),
				.m_axi4_awprot		(axi4_mem0_awprot),
				.m_axi4_awqos		(axi4_mem0_awqos),
				.m_axi4_awregion	(),
				.m_axi4_awsize		(axi4_mem0_awsize),
				.m_axi4_awvalid		(axi4_mem0_awvalid),
				.m_axi4_awready		(axi4_mem0_awready),
				.m_axi4_wstrb		(axi4_mem0_wstrb),
				.m_axi4_wdata		(axi4_mem0_wdata),
				.m_axi4_wlast		(axi4_mem0_wlast),
				.m_axi4_wvalid		(axi4_mem0_wvalid),
				.m_axi4_wready		(axi4_mem0_wready),
				.m_axi4_bid			(axi4_mem0_bid),
				.m_axi4_bresp		(axi4_mem0_bresp),
				.m_axi4_bvalid		(axi4_mem0_bvalid),
				.m_axi4_bready		(axi4_mem0_bready),
				
				/*
				.s_axi4s_aresetn	(axi4s_cam_aresetn),
				.s_axi4s_aclk		(axi4s_cam_aclk),
				.s_axi4s_tuser		(axi4s_rgb_tuser),
				.s_axi4s_tlast		(axi4s_rgb_tlast),
				.s_axi4s_tdata		({
										axi4s_rgb_tdata[39:32],
										axi4s_rgb_tdata[29:22],
										axi4s_rgb_tdata[19:12],
										axi4s_rgb_tdata[ 9: 2]
									}),
				.s_axi4s_tvalid		(axi4s_rgb_tvalid),
				.s_axi4s_tready		(axi4s_rgb_tready),
				*/
				
				.s_axi4s_aresetn	(axi4s_cam_aresetn),
				.s_axi4s_aclk		(axi4s_cam_aclk),
				.s_axi4s_tuser		(axi4s_int_tuser),
				.s_axi4s_tlast		(axi4s_int_tlast),
				.s_axi4s_tdata		({8'd0, axi4s_int_tdata}),
				.s_axi4s_tvalid		(axi4s_int_tvalid),
				.s_axi4s_tready		(axi4s_int_tready), // (axi4s_rgb_tready),
				
				
				.s_wb_rst_i			(wb_rst_o),
				.s_wb_clk_i			(wb_clk_o),
				.s_wb_adr_i			(wb_host_adr_o[7:0]),
				.s_wb_dat_o			(wb_vdmaw_dat_o),
				.s_wb_dat_i			(wb_host_dat_o),
				.s_wb_we_i			(wb_host_we_o),
				.s_wb_sel_i			(wb_host_sel_o),
				.s_wb_stb_i			(wb_vdmaw_stb_i),
				.s_wb_ack_o			(wb_vdmaw_ack_o),
				.out_irq			(),
				
				.trig_reset			(wb_rst_o),
				.trig_clk			(wb_clk_o),
				.trig_start			()
			);
	
	
	
	// ----------------------------------------
	//  VOUT
	// ----------------------------------------
	
	localparam	VOUT_X_NUM = 1280;
	localparam	VOUT_Y_NUM = 720;
	
	
	wire	[31:0]					axi4s_vout_tdata;
	wire							axi4s_vout_tlast;
	wire	[0:0]					axi4s_vout_tuser;
	wire							axi4s_vout_tvalid;
	wire							axi4s_vout_tready;
	
	/*
	jelly_pattern_generator_axi4s
			#(
				.AXI4S_DATA_WIDTH	(24),
				.X_NUM				(VOUT_X_NUM),
				.Y_NUM				(VOUT_Y_NUM),
				.X_WIDTH			(12),
				.Y_WIDTH			(12)
			)
		i_pattern_generator_axi4s
			(
				.aresetn			(~vout_reset),
				.aclk				(vout_clk),
				
				.enable				(1'b1),
				.busy				(),
				
				.m_axi4s_tdata		(axi4s_vout_tdata),
				.m_axi4s_tlast		(axi4s_vout_tlast),
				.m_axi4s_tuser		(axi4s_vout_tuser),
				.m_axi4s_tvalid		(axi4s_vout_tvalid),
				.m_axi4s_tready		(axi4s_vout_tready)
			);
	*/
	
	
	// DMA read
	wire	[31:0]			wb_vdmar_dat_o;
	wire					wb_vdmar_stb_i;
	wire					wb_vdmar_ack_o;
	
	jelly_vdma_axi4_to_axi4s
			#(
				.ASYNC				(1),
				.FIFO_PTR_WIDTH 	(9),
				
				.PIXEL_SIZE 		(2),	// 0:8bit, 1:16bit, 2:32bit, 3:64bit ...
				
				.AXI4_ID_WIDTH		(6),
				.AXI4_ADDR_WIDTH	(32),
				.AXI4_DATA_SIZE 	(3),	// 0:8bit, 1:16bit, 2:32bit, 3:64bit ...
				
				.AXI4S_DATA_SIZE	(2),	// 0:8bit, 1:16bit, 2:32bit, 3:64bit ...
				.AXI4S_USER_WIDTH	(1),
				
				.AXI4_AR_REGS		(1),
				.AXI4_R_REGS		(1),
				.AXI4S_REGS 		(1),
				
				.INDEX_WIDTH		(8),
				.STRIDE_WIDTH		(16),
				.H_WIDTH			(14),
				.V_WIDTH			(14),
				
				.WB_ADR_WIDTH		(8),
				.WB_DAT_WIDTH		(32),
				
				.TRIG_ASYNC 		(1),	// WISHBONE�Ɣ񓯊��̏ꍇ
				.TRIG_START_ENABLE	(0),
				
				.INIT_CTL_CONTROL	(4'b0000),
				.INIT_PARAM_ADDR	(32'h3000_0000),
				.INIT_PARAM_STRIDE	(8192),
				.INIT_PARAM_WIDTH	(VOUT_X_NUM),
				.INIT_PARAM_HEIGHT	(VOUT_Y_NUM),
				.INIT_PARAM_ARLEN	(8'h07)
			)
		i_vdma_axi4_to_axi4s
			(
				.m_axi4_aresetn		(axi4_mem_aresetn),
				.m_axi4_aclk		(axi4_mem_aclk),
				.m_axi4_arid		(axi4_mem0_arid),
				.m_axi4_araddr		(axi4_mem0_araddr),
				.m_axi4_arlen		(axi4_mem0_arlen),
				.m_axi4_arsize		(axi4_mem0_arsize),
				.m_axi4_arburst		(axi4_mem0_arburst),
				.m_axi4_arlock		(axi4_mem0_arlock),
				.m_axi4_arcache		(axi4_mem0_arcache),
				.m_axi4_arprot		(axi4_mem0_arprot),
				.m_axi4_arqos		(axi4_mem0_arqos),
				.m_axi4_arregion	(axi4_mem0_arregion),
				.m_axi4_arvalid		(axi4_mem0_arvalid),
				.m_axi4_arready		(axi4_mem0_arready),
				.m_axi4_rid			(axi4_mem0_rid),
				.m_axi4_rdata		(axi4_mem0_rdata),
				.m_axi4_rresp		(axi4_mem0_rresp),
				.m_axi4_rlast		(axi4_mem0_rlast),
				.m_axi4_rvalid		(axi4_mem0_rvalid),
				.m_axi4_rready		(axi4_mem0_rready),
				
				.m_axi4s_aresetn	(~vout_reset),
				.m_axi4s_aclk		(vout_clk),
				.m_axi4s_tdata		(axi4s_vout_tdata),
				.m_axi4s_tlast		(axi4s_vout_tlast),
				.m_axi4s_tuser		(axi4s_vout_tuser),
				.m_axi4s_tvalid		(axi4s_vout_tvalid),
				.m_axi4s_tready		(axi4s_vout_tready),
				
				.s_wb_rst_i			(wb_rst_o),
				.s_wb_clk_i			(wb_clk_o),
				.s_wb_adr_i			(wb_host_adr_o[7:0]),
				.s_wb_dat_i			(wb_host_dat_o),
				.s_wb_dat_o			(wb_vdmar_dat_o),
				.s_wb_we_i			(wb_host_we_o),
				.s_wb_sel_i			(wb_host_sel_o),
				.s_wb_stb_i			(wb_vdmar_stb_i),
				.s_wb_ack_o			(wb_vdmar_ack_o),
				.out_irq			(),
				
				.trig_reset			(wb_rst_o),
				.trig_clk			(wb_clk_o),
				.trig_start			(0)
			);
	
	
//	// read �͖��g�p
//	assign axi4_mem0_arid     = 0;
//	assign axi4_mem0_araddr   = 0;
//	assign axi4_mem0_arburst  = 0;
//	assign axi4_mem0_arcache  = 0;
//	assign axi4_mem0_arlen    = 0;
//	assign axi4_mem0_arlock   = 0;
//	assign axi4_mem0_arprot   = 0;
//	assign axi4_mem0_arqos    = 0;
//	assign axi4_mem0_arregion = 0;
//	assign axi4_mem0_arsize   = 0;
//	assign axi4_mem0_arvalid  = 0;
//	assign axi4_mem0_rready   = 0;
	
	
	wire					vout_vsgen_vsync;
	wire					vout_vsgen_hsync;
	wire					vout_vsgen_de;
	
	wire	[31:0]			wb_vsgen_dat_o;
	wire					wb_vsgen_stb_i;
	wire					wb_vsgen_ack_o;
	
	jelly_vsync_generator
			#(
				.WB_ADR_WIDTH		(8),
				.WB_DAT_WIDTH		(32),
				.INIT_CTL_CONTROL	(1'b0),
				
				.INIT_HTOTAL		(1650),
				.INIT_HDISP_START	(0),
				.INIT_HDISP_END		(VOUT_X_NUM),
				.INIT_HSYNC_START	(1390),
				.INIT_HSYNC_END		(1430),
				.INIT_HSYNC_POL		(1),
				.INIT_VTOTAL		(750),
				.INIT_VDISP_START	(0),
				.INIT_VDISP_END		(VOUT_Y_NUM),
				.INIT_VSYNC_START	(725),
				.INIT_VSYNC_END		(730),
				.INIT_VSYNC_POL		(1)
			)
		i_vsync_generator
			(
				.reset				(vout_reset),
				.clk				(vout_clk),
				
				.out_vsync			(vout_vsgen_vsync),
				.out_hsync			(vout_vsgen_hsync),
				.out_de				(vout_vsgen_de),
				
				.s_wb_rst_i			(wb_rst_o),
				.s_wb_clk_i			(wb_clk_o),
				.s_wb_adr_i			(wb_host_adr_o[7:0]),
				.s_wb_dat_o			(wb_vsgen_dat_o),
				.s_wb_dat_i			(wb_host_dat_o),
				.s_wb_we_i			(wb_host_we_o),
				.s_wb_sel_i			(wb_host_sel_o),
				.s_wb_stb_i			(wb_vsgen_stb_i),
				.s_wb_ack_o			(wb_vsgen_ack_o)
			);
	
	
	(* MARK_DEBUG="true" *)	wire			vout_vsync;
	(* MARK_DEBUG="true" *)	wire			vout_hsync;
	(* MARK_DEBUG="true" *)	wire			vout_de;
	(* MARK_DEBUG="true" *)	wire	[23:0]	vout_data;
	(* MARK_DEBUG="true" *)	wire	[3:0]	vout_ctl;
	
	jelly_vout_axi4s
			#(
				.WIDTH				(24)
			)
		i_vout_axi4s
			(
				.reset				(vout_reset),
				.clk				(vout_clk),
				
				.s_axi4s_tuser		(axi4s_vout_tuser),
				.s_axi4s_tlast		(axi4s_vout_tlast),
				.s_axi4s_tdata		(axi4s_vout_tdata[23:0]),
				.s_axi4s_tvalid		(axi4s_vout_tvalid),
				.s_axi4s_tready		(axi4s_vout_tready),
				
				.in_vsync			(vout_vsgen_vsync),
				.in_hsync			(vout_vsgen_hsync),
				.in_de				(vout_vsgen_de),
				.in_ctl				(4'd0),
				
				.out_vsync			(vout_vsync),
				.out_hsync			(vout_hsync),
				.out_de				(vout_de),
				.out_data			(vout_data),
				.out_ctl			(vout_ctl)
			);
	
	jelly_dvi_tx
		i_dvi_tx
			(
				.reset				(vout_reset),
				.clk				(vout_clk),
				.clk_x5				(vout_clk_x5),
				
				.in_vsync			(vout_vsync),
				.in_hsync			(vout_hsync),
				.in_de				(vout_de),
				.in_data			(vout_data),
				.in_ctl				(4'd0),
				
				.out_clk_p			(hdmi_tx_clk_p),
				.out_clk_n			(hdmi_tx_clk_n),
				.out_data_p			(hdmi_tx_data_p),
				.out_data_n			(hdmi_tx_data_n)
			);
	
	
	// ----------------------------------------
	//  �P���_���v
	// ----------------------------------------
	/*
	// FIFO
	(* MARK_DEBUG = "true" *)	wire	[7:0]		fifo_dl0_rxdatahs;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl0_rxvalidhs;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl0_rxactivehs;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl0_rxsynchs;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl0_errsoths;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl0_errsotsynchs;
	(* MARK_DEBUG = "true" *)	wire	[7:0]		fifo_dl1_rxdatahs;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl1_rxvalidhs;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl1_rxactivehs;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl1_rxsynchs;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl1_errsoths;
	(* MARK_DEBUG = "true" *)	wire				fifo_dl1_errsotsynchs;
	(* MARK_DEBUG = "true" *)	wire				fifo_valid;
	
	jelly_fifo_async_fwtf
			#(
				.DATA_WIDTH			((5+8)*2),
				.PTR_WIDTH			(6),
				.DOUT_REGS			(0),
				.RAM_TYPE			("distributed"),
				.SLAVE_REGS			(0),
				.MASTER_REGS		(1)
			)
		i_fifo_async_fwtf
			(
				.s_reset			(dphy_reset),
				.s_clk				(dphy_clk),
				.s_data				({
										dl0_rxdatahs,
										dl0_rxvalidhs,
										dl0_rxactivehs,
										dl0_rxsynchs,
										dl0_errsoths,
										dl0_errsotsynchs,
										dl1_rxdatahs,
										dl1_rxvalidhs,
										dl1_rxactivehs,
										dl1_rxsynchs,
										dl1_errsoths,
										dl1_errsotsynchs
									}),
				.s_valid			(1'b1),
				.s_ready			(),
				.s_free_count		(),
				
				.m_reset			(~axi4_mem_aresetn),
				.m_clk				(axi4_mem_aclk),
				.m_data				({
										fifo_dl0_rxdatahs,
										fifo_dl0_rxvalidhs,
										fifo_dl0_rxactivehs,
										fifo_dl0_rxsynchs,
										fifo_dl0_errsoths,
										fifo_dl0_errsotsynchs,
										fifo_dl1_rxdatahs,
										fifo_dl1_rxvalidhs,
										fifo_dl1_rxactivehs,
										fifo_dl1_rxsynchs,
										fifo_dl1_errsoths,
										fifo_dl1_errsotsynchs
									}),
				.m_valid			(fifo_valid),
				.m_ready			(1'b1),
				.m_data_count		()
			);
	
	
	(* MARK_DEBUG = "true" *)	wire	[0:0]			axi4s_memw_tuser;
	(* MARK_DEBUG = "true" *)	wire					axi4s_memw_tlast;
	(* MARK_DEBUG = "true" *)	wire	[31:0]			axi4s_memw_tdata;
	(* MARK_DEBUG = "true" *)	wire					axi4s_memw_tvalid;
	(* MARK_DEBUG = "true" *)	wire					axi4s_memw_tready;
	
	assign axi4s_memw_tuser       = fifo_dl0_rxsynchs;
	assign axi4s_memw_tlast       = 1'b0;
	assign axi4s_memw_tdata[15:0] = {
										fifo_dl0_errsotsynchs,
										fifo_dl0_errsoths,
										fifo_dl0_rxsynchs,
										fifo_dl0_rxactivehs,
										fifo_dl0_rxvalidhs,
										fifo_dl0_rxdatahs
									};
	assign axi4s_memw_tdata[31:16] = {
										fifo_dl1_errsotsynchs,
										fifo_dl1_errsoths,
										fifo_dl1_rxsynchs,
										fifo_dl1_rxactivehs,
										fifo_dl1_rxvalidhs,
										fifo_dl1_rxdatahs
									};
	
	assign axi4s_memw_tvalid       = fifo_valid;
	
	
	
	(* MARK_DEBUG = "true" *)	wire	[31:0]			wb_vdmaw_dat_o;
	(* MARK_DEBUG = "true" *)	wire					wb_vdmaw_stb_i;
	(* MARK_DEBUG = "true" *)	wire					wb_vdmaw_ack_o;
	
	reg				vdmaw_enable;
	wire			vdmaw_busy;
	
	always @(posedge wb_clk_o ) begin
		if ( wb_rst_o ) begin
			vdmaw_enable <= 0;
		end
		else begin
			vdmaw_enable <= 0;
			if ( wb_vdmaw_stb_i && wb_host_we_o ) begin
				vdmaw_enable <= wb_host_dat_o;
			end
		end
	end
	
	assign wb_vdmaw_dat_o = vdmaw_busy;
	assign wb_vdmaw_ack_o = wb_vdmaw_stb_i;
	
	reg				vdmaw_enable_ff0, vdmaw_enable_ff1;
	always @(posedge axi4_mem_aclk) begin
		vdmaw_enable_ff0 <= vdmaw_enable;
		vdmaw_enable_ff1 <= vdmaw_enable_ff0;
	end
	
	
	jelly_axi4_dma_writer
			#(
				.AXI4_ID_WIDTH		(6),
				.AXI4_ADDR_WIDTH	(32),
				.AXI4_DATA_SIZE		(3)		// 0:8bit, 1:16bit, 2:32bit ...
			)
		i_axi4_dma_writer
			(
				.aresetn			(axi4_mem_aresetn),
				.aclk				(axi4_mem_aclk),
				
				.enable				(vdmaw_enable_ff1),
				.busy				(vdmaw_busy),
				
				.queue_counter		(0),
				
				.param_addr			(32'h1000_0000),
				.param_count		(64*1024*1024),
				.param_maxlen		(7),
				.param_wstrb		(8'hff),
				
				.m_axi4_awid		(axi4_mem0_awid),
				.m_axi4_awaddr		(axi4_mem0_awaddr),
				.m_axi4_awburst		(axi4_mem0_awburst),
				.m_axi4_awcache		(axi4_mem0_awcache),
				.m_axi4_awlen		(axi4_mem0_awlen),
				.m_axi4_awlock		(axi4_mem0_awlock),
				.m_axi4_awprot		(axi4_mem0_awprot),
				.m_axi4_awqos		(axi4_mem0_awqos),
				.m_axi4_awregion	(),
				.m_axi4_awsize		(axi4_mem0_awsize),
				.m_axi4_awvalid		(axi4_mem0_awvalid),
				.m_axi4_awready		(axi4_mem0_awready),
				.m_axi4_wstrb		(axi4_mem0_wstrb),
				.m_axi4_wdata		(axi4_mem0_wdata),
				.m_axi4_wlast		(axi4_mem0_wlast),
				.m_axi4_wvalid		(axi4_mem0_wvalid),
				.m_axi4_wready		(axi4_mem0_wready),
				.m_axi4_bid			(axi4_mem0_bid),
				.m_axi4_bresp		(axi4_mem0_bresp),
				.m_axi4_bvalid		(axi4_mem0_bvalid),
				.m_axi4_bready		(axi4_mem0_bready),
				
				.s_axi4s_tdata		({32'd0, axi4s_memw_tdata}),
				.s_axi4s_tvalid		(axi4s_memw_tvalid),
				.s_axi4s_tready		(axi4s_memw_tready)
			);
	*/
	
	
	
	

	
	
	
	// ----------------------------------------
	//  WISHBONE address decoder
	// ----------------------------------------
	
	assign wb_gid_stb_i   = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4000_0);
	assign wb_vdmaw_stb_i = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4001_0);
	assign wb_norm_stb_i  = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4001_1);
	assign wb_rgb_stb_i   = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4001_2);
	assign wb_mnist_stb_i = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4001_8);
	assign wb_mcol_stb_i  = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4001_9);
	assign wb_int_stb_i   = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4001_a);
	assign wb_vdmar_stb_i = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4002_0);
	assign wb_vsgen_stb_i = wb_host_stb_o & (wb_host_adr_o[29:10] == 20'h4002_1);
	
	
	assign wb_host_dat_i  = wb_gid_stb_i   ? wb_gid_dat_o   :
	                        wb_vdmaw_stb_i ? wb_vdmaw_dat_o :
	                        wb_norm_stb_i  ? wb_norm_dat_o  :
	                        wb_rgb_stb_i   ? wb_rgb_dat_o   :
	                        wb_mnist_stb_i ? wb_mnist_dat_o :
	                        wb_mcol_stb_i  ? wb_mcol_dat_o  :
	                        wb_int_stb_i   ? wb_int_dat_o   :
	                        wb_vdmar_stb_i ? wb_vdmar_dat_o :
	                        wb_vsgen_stb_i ? wb_vsgen_dat_o :
	                        32'h0000_0000;
	
	assign wb_host_ack_i  = wb_gid_stb_i   ? wb_gid_ack_o   :
	                        wb_vdmaw_stb_i ? wb_vdmaw_ack_o :
	                        wb_norm_stb_i  ? wb_norm_ack_o  :
	                        wb_rgb_stb_i   ? wb_rgb_ack_o   :
	                        wb_mnist_stb_i ? wb_mnist_ack_o :
	                        wb_mcol_stb_i  ? wb_mcol_ack_o  :
	                        wb_int_stb_i   ? wb_int_ack_o   :
	                        wb_vdmar_stb_i ? wb_vdmar_ack_o :
	                        wb_vsgen_stb_i ? wb_vsgen_ack_o :
	                        wb_host_stb_o;
	
	
	
	// ----------------------------------------
	//  Debug
	// ----------------------------------------
	
	reg		[31:0]		reg_counter_rxbyteclkhs;
	always @(posedge rxbyteclkhs)	reg_counter_rxbyteclkhs <= reg_counter_rxbyteclkhs + 1;
	
	reg		[31:0]		reg_counter_clk200;
	always @(posedge sys_clk200)	reg_counter_clk200 <= reg_counter_clk200 + 1;
	
	reg		[31:0]		reg_counter_clk100;
	always @(posedge sys_clk100)	reg_counter_clk100 <= reg_counter_clk100 + 1;
	
	
	reg		frame_toggle = 0;
	always @(posedge axi4s_cam_aclk) begin
		if ( axi4s_csi2_tuser[0] && axi4s_csi2_tvalid && axi4s_csi2_tready ) begin
			frame_toggle <= ~frame_toggle;
		end
	end
	
	
	assign led[0] = reg_counter_rxbyteclkhs[24];
	assign led[1] = reg_counter_clk200[24];
	assign led[2] = reg_counter_clk100[24];
	assign led[3] = frame_toggle;
	
	assign pmod_a[0]   = frame_toggle;
	assign pmod_a[1]   = reg_counter_rxbyteclkhs[5];
	assign pmod_a[2]   = reg_counter_clk200[5];
	assign pmod_a[3]   = reg_counter_clk100[5];
	assign pmod_a[7:4] = 0;
	
	
	(* MARK_DEBUG = "true" *) reg	dbg_clk200;
	(* MARK_DEBUG = "true" *) reg	dbg_clk100;
	(* MARK_DEBUG = "true" *) reg	dbg_rxbyteclkhs;
	always @(posedge sys_clk100) begin
		dbg_clk200       <= reg_counter_clk200[5];
		dbg_clk100       <= reg_counter_clk100[5];
		dbg_rxbyteclkhs  <= reg_counter_rxbyteclkhs[5];
	end
	
	
endmodule


`default_nettype wire

