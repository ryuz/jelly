

module OSER10
    (
        output  wire    Q    ,
        input   wire    D0   ,
        input   wire    D1   ,
        input   wire    D2   ,
        input   wire    D3   ,
        input   wire    D4   ,
        input   wire    D5   ,
        input   wire    D6   ,
        input   wire    D7   ,
        input   wire    D8   ,
        input   wire    D9   ,
        input   wire    PCLK ,
        input   wire    FCLK ,
        input   wire    RESET
    );

endmodule
