// ---------------------------------------------------------------------------
//  Jelly  -- the soft-core processor system
//   image processing
//
//                                 Copyright (C) 2008-2016 by Ryuji Fuchikami
//                                 http://ryuz.my.coocan.jp/
// ---------------------------------------------------------------------------



`timescale 1ns / 1ps
`default_nettype none


module jelly_img_demosaic_acpi_rb_core
		#(
			parameter	USER_WIDTH = 0,
			parameter	DATA_WIDTH = 10,
			parameter	MAX_X_NUM  = 4096,
			parameter	USE_VALID  = 0,
			
			parameter	USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
		)
		(
			input	wire							reset,
			input	wire							clk,
			input	wire							cke,
			
			input	wire	[1:0]					param_phase,
			
			input	wire							s_img_line_first,
			input	wire							s_img_line_last,
			input	wire							s_img_pixel_first,
			input	wire							s_img_pixel_last,
			input	wire							s_img_de,
			input	wire	[USER_BITS-1:0]			s_img_user,
			input	wire	[DATA_WIDTH-1:0]		s_img_raw,
			input	wire	[DATA_WIDTH-1:0]		s_img_g,
			input	wire							s_img_valid,
			
			output	wire							m_img_line_first,
			output	wire							m_img_line_last,
			output	wire							m_img_pixel_first,
			output	wire							m_img_pixel_last,
			output	wire							m_img_de,
			output	wire	[USER_BITS-1:0]			m_img_user,
			output	wire	[DATA_WIDTH-1:0]		m_img_raw,
			output	wire	[DATA_WIDTH-1:0]		m_img_r,
			output	wire	[DATA_WIDTH-1:0]		m_img_g,
			output	wire	[DATA_WIDTH-1:0]		m_img_b,
			output	wire							m_img_valid
		);
	
	
	wire							img_blk_line_first;
	wire							img_blk_line_last;
	wire							img_blk_pixel_first;
	wire							img_blk_pixel_last;
	wire	[USER_BITS-1:0]			img_blk_user;
	wire							img_blk_de;
	wire	[3*3*2*DATA_WIDTH-1:0]	img_blk_data;
	wire							img_blk_valid;
	
	jelly_img_blk_buffer
			#(
				.DATA_WIDTH			(2*DATA_WIDTH),
				.LINE_NUM			(3),
				.PIXEL_NUM			(3),
				.MAX_X_NUM			(MAX_X_NUM),
				.RAM_TYPE			("block"),
				.BORDER_MODE		("REFLECT_101")
			)
		i_img_blk_buffer
			(
				.reset				(reset),
				.clk				(clk),
				.cke				(cke),
				
				.s_img_line_first	(s_img_line_first),
				.s_img_line_last	(s_img_line_last),
				.s_img_pixel_first	(s_img_pixel_first),
				.s_img_pixel_last	(s_img_pixel_last),
				.s_img_de			(s_img_de),
				.s_img_user			(s_img_user),
				.s_img_data			({s_img_g, s_img_raw}),
				.s_img_valid		(s_img_valid),
				
				.m_img_line_first	(img_blk_line_first),
				.m_img_line_last	(img_blk_line_last),
				.m_img_pixel_first	(img_blk_pixel_first),
				.m_img_pixel_last	(img_blk_pixel_last),
				.m_img_de			(img_blk_de),
				.m_img_user			(img_blk_user),
				.m_img_data			(img_blk_data),
				.m_img_valid		(img_blk_valid)
			);
	
	
	jelly_img_demosaic_acpi_rb_unit
			#(
				.DATA_WIDTH			(DATA_WIDTH)
			)
		i_img_demosaic_acpi_rb_unit
			(
				.reset				(reset),
				.clk				(clk),
				.cke				(cke),
				
				.param_phase		(param_phase),
				
				.in_line_first		(img_blk_line_first  & img_blk_valid),
				.in_pixel_first		(img_blk_pixel_first & img_blk_valid),
				.in_data			(img_blk_data),
				
				.out_raw			(m_img_raw),
				.out_r				(m_img_r),
				.out_g				(m_img_g),
				.out_b				(m_img_b)
			);
	
	jelly_img_delay
			#(
				.USER_WIDTH			(USER_WIDTH),
				.LATENCY			(6),
				.USE_VALID			(USE_VALID)
			)
		i_img_delay
			(
				.reset				(reset),
				.clk				(clk),
				.cke				(cke),
				
				.s_img_line_first	(img_blk_line_first),
				.s_img_line_last	(img_blk_line_last),
				.s_img_pixel_first	(img_blk_pixel_first),
				.s_img_pixel_last	(img_blk_pixel_last),
				.s_img_de			(img_blk_de),
				.s_img_user			(img_blk_user),
				.s_img_valid		(img_blk_valid),
				
				.m_img_line_first	(m_img_line_first),
				.m_img_line_last	(m_img_line_last),
				.m_img_pixel_first	(m_img_pixel_first),
				.m_img_pixel_last	(m_img_pixel_last),
				.m_img_de			(m_img_de),
				.m_img_user			(m_img_user),
				.m_img_valid		(m_img_valid)
			);
	
	
endmodule


`default_nettype wire


// end of file
