
`timescale 1ns / 1ps
`default_nettype none

module clk_wiz_0
        (
            input   var logic clk_in1,
            output  var logic clk_out1,
            output  var logic clk_out2,
            output  var logic clk_out3
        );


endmodule

`default_nettype wire

// end of file
