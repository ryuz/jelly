// ---------------------------------------------------------------------------
//  Jelly  -- The platform for real-time computing
//
//                                 Copyright (C) 2008-2020 by Ryuji Fuchikami
//                                 https://github.com/ryuz/jelly.git
// ---------------------------------------------------------------------------



`timescale 1ns / 1ps
`default_nettype none


// colormap
module jelly_colormap_table
        #(
            parameter   COLORMAP = "JET"   // "HSV"
        )
        (
            input   wire    [7:0]       in_data,
            output  reg     [23:0]      out_data
        );
    
    always @* begin
        if ( COLORMAP == "HSV" ) begin
            case ( in_data )
            8'h00:  out_data = 24'h00_00_ff;
            8'h01:  out_data = 24'h00_06_ff;
            8'h02:  out_data = 24'h00_0c_ff;
            8'h03:  out_data = 24'h00_12_ff;
            8'h04:  out_data = 24'h00_18_ff;
            8'h05:  out_data = 24'h00_1e_ff;
            8'h06:  out_data = 24'h00_24_ff;
            8'h07:  out_data = 24'h00_2a_ff;
            8'h08:  out_data = 24'h00_30_ff;
            8'h09:  out_data = 24'h00_36_ff;
            8'h0a:  out_data = 24'h00_3c_ff;
            8'h0b:  out_data = 24'h00_42_ff;
            8'h0c:  out_data = 24'h00_48_ff;
            8'h0d:  out_data = 24'h00_4e_ff;
            8'h0e:  out_data = 24'h00_54_ff;
            8'h0f:  out_data = 24'h00_5a_ff;
            8'h10:  out_data = 24'h00_60_ff;
            8'h11:  out_data = 24'h00_66_ff;
            8'h12:  out_data = 24'h00_6c_ff;
            8'h13:  out_data = 24'h00_72_ff;
            8'h14:  out_data = 24'h00_78_ff;
            8'h15:  out_data = 24'h00_7e_ff;
            8'h16:  out_data = 24'h00_84_ff;
            8'h17:  out_data = 24'h00_8a_ff;
            8'h18:  out_data = 24'h00_90_ff;
            8'h19:  out_data = 24'h00_96_ff;
            8'h1a:  out_data = 24'h00_9c_ff;
            8'h1b:  out_data = 24'h00_a2_ff;
            8'h1c:  out_data = 24'h00_a8_ff;
            8'h1d:  out_data = 24'h00_ae_ff;
            8'h1e:  out_data = 24'h00_b4_ff;
            8'h1f:  out_data = 24'h00_ba_ff;
            8'h20:  out_data = 24'h00_c0_ff;
            8'h21:  out_data = 24'h00_c6_ff;
            8'h22:  out_data = 24'h00_cc_ff;
            8'h23:  out_data = 24'h00_d2_ff;
            8'h24:  out_data = 24'h00_d8_ff;
            8'h25:  out_data = 24'h00_de_ff;
            8'h26:  out_data = 24'h00_e4_ff;
            8'h27:  out_data = 24'h00_ea_ff;
            8'h28:  out_data = 24'h00_f0_ff;
            8'h29:  out_data = 24'h00_f4_fd;
            8'h2a:  out_data = 24'h00_f7_fa;
            8'h2b:  out_data = 24'h00_fa_f7;
            8'h2c:  out_data = 24'h00_fd_f4;
            8'h2d:  out_data = 24'h00_ff_f0;
            8'h2e:  out_data = 24'h00_ff_ea;
            8'h2f:  out_data = 24'h00_ff_e4;
            8'h30:  out_data = 24'h00_ff_de;
            8'h31:  out_data = 24'h00_ff_d8;
            8'h32:  out_data = 24'h00_ff_d2;
            8'h33:  out_data = 24'h00_ff_cc;
            8'h34:  out_data = 24'h00_ff_c6;
            8'h35:  out_data = 24'h00_ff_c0;
            8'h36:  out_data = 24'h00_ff_ba;
            8'h37:  out_data = 24'h00_ff_b4;
            8'h38:  out_data = 24'h00_ff_ae;
            8'h39:  out_data = 24'h00_ff_a8;
            8'h3a:  out_data = 24'h00_ff_a2;
            8'h3b:  out_data = 24'h00_ff_9c;
            8'h3c:  out_data = 24'h00_ff_96;
            8'h3d:  out_data = 24'h00_ff_90;
            8'h3e:  out_data = 24'h00_ff_8a;
            8'h3f:  out_data = 24'h00_ff_84;
            8'h40:  out_data = 24'h00_ff_7e;
            8'h41:  out_data = 24'h00_ff_78;
            8'h42:  out_data = 24'h00_ff_72;
            8'h43:  out_data = 24'h00_ff_6c;
            8'h44:  out_data = 24'h00_ff_66;
            8'h45:  out_data = 24'h00_ff_60;
            8'h46:  out_data = 24'h00_ff_5a;
            8'h47:  out_data = 24'h00_ff_54;
            8'h48:  out_data = 24'h00_ff_4e;
            8'h49:  out_data = 24'h00_ff_48;
            8'h4a:  out_data = 24'h00_ff_42;
            8'h4b:  out_data = 24'h00_ff_3c;
            8'h4c:  out_data = 24'h00_ff_36;
            8'h4d:  out_data = 24'h00_ff_30;
            8'h4e:  out_data = 24'h00_ff_2a;
            8'h4f:  out_data = 24'h00_ff_24;
            8'h50:  out_data = 24'h00_ff_1e;
            8'h51:  out_data = 24'h00_ff_18;
            8'h52:  out_data = 24'h00_ff_12;
            8'h53:  out_data = 24'h00_ff_0c;
            8'h54:  out_data = 24'h00_ff_06;
            8'h55:  out_data = 24'h00_ff_00;
            8'h56:  out_data = 24'h06_ff_00;
            8'h57:  out_data = 24'h0c_ff_00;
            8'h58:  out_data = 24'h12_ff_00;
            8'h59:  out_data = 24'h18_ff_00;
            8'h5a:  out_data = 24'h1e_ff_00;
            8'h5b:  out_data = 24'h24_ff_00;
            8'h5c:  out_data = 24'h2a_ff_00;
            8'h5d:  out_data = 24'h30_ff_00;
            8'h5e:  out_data = 24'h36_ff_00;
            8'h5f:  out_data = 24'h3c_ff_00;
            8'h60:  out_data = 24'h42_ff_00;
            8'h61:  out_data = 24'h48_ff_00;
            8'h62:  out_data = 24'h4e_ff_00;
            8'h63:  out_data = 24'h54_ff_00;
            8'h64:  out_data = 24'h5a_ff_00;
            8'h65:  out_data = 24'h60_ff_00;
            8'h66:  out_data = 24'h66_ff_00;
            8'h67:  out_data = 24'h6c_ff_00;
            8'h68:  out_data = 24'h72_ff_00;
            8'h69:  out_data = 24'h78_ff_00;
            8'h6a:  out_data = 24'h7e_ff_00;
            8'h6b:  out_data = 24'h84_ff_00;
            8'h6c:  out_data = 24'h8a_ff_00;
            8'h6d:  out_data = 24'h90_ff_00;
            8'h6e:  out_data = 24'h96_ff_00;
            8'h6f:  out_data = 24'h9c_ff_00;
            8'h70:  out_data = 24'ha2_ff_00;
            8'h71:  out_data = 24'ha8_ff_00;
            8'h72:  out_data = 24'hae_ff_00;
            8'h73:  out_data = 24'hb4_ff_00;
            8'h74:  out_data = 24'hba_ff_00;
            8'h75:  out_data = 24'hc0_ff_00;
            8'h76:  out_data = 24'hc6_ff_00;
            8'h77:  out_data = 24'hcc_ff_00;
            8'h78:  out_data = 24'hd2_ff_00;
            8'h79:  out_data = 24'hd8_ff_00;
            8'h7a:  out_data = 24'hde_ff_00;
            8'h7b:  out_data = 24'he4_ff_00;
            8'h7c:  out_data = 24'hea_ff_00;
            8'h7d:  out_data = 24'hf0_ff_00;
            8'h7e:  out_data = 24'hf4_fd_00;
            8'h7f:  out_data = 24'hf7_fa_00;
            8'h80:  out_data = 24'hfa_f7_00;
            8'h81:  out_data = 24'hfd_f4_00;
            8'h82:  out_data = 24'hff_f0_00;
            8'h83:  out_data = 24'hff_ea_00;
            8'h84:  out_data = 24'hff_e4_00;
            8'h85:  out_data = 24'hff_de_00;
            8'h86:  out_data = 24'hff_d8_00;
            8'h87:  out_data = 24'hff_d2_00;
            8'h88:  out_data = 24'hff_cc_00;
            8'h89:  out_data = 24'hff_c6_00;
            8'h8a:  out_data = 24'hff_c0_00;
            8'h8b:  out_data = 24'hff_ba_00;
            8'h8c:  out_data = 24'hff_b4_00;
            8'h8d:  out_data = 24'hff_ae_00;
            8'h8e:  out_data = 24'hff_a8_00;
            8'h8f:  out_data = 24'hff_a2_00;
            8'h90:  out_data = 24'hff_9c_00;
            8'h91:  out_data = 24'hff_96_00;
            8'h92:  out_data = 24'hff_90_00;
            8'h93:  out_data = 24'hff_8a_00;
            8'h94:  out_data = 24'hff_84_00;
            8'h95:  out_data = 24'hff_7e_00;
            8'h96:  out_data = 24'hff_78_00;
            8'h97:  out_data = 24'hff_72_00;
            8'h98:  out_data = 24'hff_6c_00;
            8'h99:  out_data = 24'hff_66_00;
            8'h9a:  out_data = 24'hff_60_00;
            8'h9b:  out_data = 24'hff_5a_00;
            8'h9c:  out_data = 24'hff_54_00;
            8'h9d:  out_data = 24'hff_4e_00;
            8'h9e:  out_data = 24'hff_48_00;
            8'h9f:  out_data = 24'hff_42_00;
            8'ha0:  out_data = 24'hff_3c_00;
            8'ha1:  out_data = 24'hff_36_00;
            8'ha2:  out_data = 24'hff_30_00;
            8'ha3:  out_data = 24'hff_2a_00;
            8'ha4:  out_data = 24'hff_24_00;
            8'ha5:  out_data = 24'hff_1e_00;
            8'ha6:  out_data = 24'hff_18_00;
            8'ha7:  out_data = 24'hff_12_00;
            8'ha8:  out_data = 24'hff_0c_00;
            8'ha9:  out_data = 24'hff_06_00;
            8'haa:  out_data = 24'hff_00_00;
            8'hab:  out_data = 24'hff_00_06;
            8'hac:  out_data = 24'hff_00_0c;
            8'had:  out_data = 24'hff_00_12;
            8'hae:  out_data = 24'hff_00_18;
            8'haf:  out_data = 24'hff_00_1e;
            8'hb0:  out_data = 24'hff_00_24;
            8'hb1:  out_data = 24'hff_00_2a;
            8'hb2:  out_data = 24'hff_00_30;
            8'hb3:  out_data = 24'hff_00_36;
            8'hb4:  out_data = 24'hff_00_3c;
            8'hb5:  out_data = 24'hff_00_42;
            8'hb6:  out_data = 24'hff_00_48;
            8'hb7:  out_data = 24'hff_00_4e;
            8'hb8:  out_data = 24'hff_00_54;
            8'hb9:  out_data = 24'hff_00_5a;
            8'hba:  out_data = 24'hff_00_60;
            8'hbb:  out_data = 24'hff_00_66;
            8'hbc:  out_data = 24'hff_00_6c;
            8'hbd:  out_data = 24'hff_00_72;
            8'hbe:  out_data = 24'hff_00_78;
            8'hbf:  out_data = 24'hff_00_7e;
            8'hc0:  out_data = 24'hff_00_84;
            8'hc1:  out_data = 24'hff_00_8a;
            8'hc2:  out_data = 24'hff_00_90;
            8'hc3:  out_data = 24'hff_00_96;
            8'hc4:  out_data = 24'hff_00_9c;
            8'hc5:  out_data = 24'hff_00_a2;
            8'hc6:  out_data = 24'hff_00_a8;
            8'hc7:  out_data = 24'hff_00_ae;
            8'hc8:  out_data = 24'hff_00_b4;
            8'hc9:  out_data = 24'hff_00_ba;
            8'hca:  out_data = 24'hff_00_c0;
            8'hcb:  out_data = 24'hff_00_c6;
            8'hcc:  out_data = 24'hff_00_cc;
            8'hcd:  out_data = 24'hff_00_d2;
            8'hce:  out_data = 24'hff_00_d8;
            8'hcf:  out_data = 24'hff_00_de;
            8'hd0:  out_data = 24'hff_00_e4;
            8'hd1:  out_data = 24'hff_00_ea;
            8'hd2:  out_data = 24'hff_00_f0;
            8'hd3:  out_data = 24'hfd_00_f4;
            8'hd4:  out_data = 24'hfa_00_f7;
            8'hd5:  out_data = 24'hf7_00_fa;
            8'hd6:  out_data = 24'hf4_00_fd;
            8'hd7:  out_data = 24'hf0_00_ff;
            8'hd8:  out_data = 24'hea_00_ff;
            8'hd9:  out_data = 24'he4_00_ff;
            8'hda:  out_data = 24'hde_00_ff;
            8'hdb:  out_data = 24'hd8_00_ff;
            8'hdc:  out_data = 24'hd2_00_ff;
            8'hdd:  out_data = 24'hcc_00_ff;
            8'hde:  out_data = 24'hc6_00_ff;
            8'hdf:  out_data = 24'hc0_00_ff;
            8'he0:  out_data = 24'hba_00_ff;
            8'he1:  out_data = 24'hb4_00_ff;
            8'he2:  out_data = 24'hae_00_ff;
            8'he3:  out_data = 24'ha8_00_ff;
            8'he4:  out_data = 24'ha2_00_ff;
            8'he5:  out_data = 24'h9c_00_ff;
            8'he6:  out_data = 24'h96_00_ff;
            8'he7:  out_data = 24'h90_00_ff;
            8'he8:  out_data = 24'h8a_00_ff;
            8'he9:  out_data = 24'h84_00_ff;
            8'hea:  out_data = 24'h7e_00_ff;
            8'heb:  out_data = 24'h78_00_ff;
            8'hec:  out_data = 24'h72_00_ff;
            8'hed:  out_data = 24'h6c_00_ff;
            8'hee:  out_data = 24'h66_00_ff;
            8'hef:  out_data = 24'h60_00_ff;
            8'hf0:  out_data = 24'h5a_00_ff;
            8'hf1:  out_data = 24'h54_00_ff;
            8'hf2:  out_data = 24'h4e_00_ff;
            8'hf3:  out_data = 24'h48_00_ff;
            8'hf4:  out_data = 24'h42_00_ff;
            8'hf5:  out_data = 24'h3c_00_ff;
            8'hf6:  out_data = 24'h36_00_ff;
            8'hf7:  out_data = 24'h30_00_ff;
            8'hf8:  out_data = 24'h2a_00_ff;
            8'hf9:  out_data = 24'h24_00_ff;
            8'hfa:  out_data = 24'h1e_00_ff;
            8'hfb:  out_data = 24'h18_00_ff;
            8'hfc:  out_data = 24'h12_00_ff;
            8'hfd:  out_data = 24'h0c_00_ff;
            8'hfe:  out_data = 24'h06_00_ff;
            8'hff:  out_data = 24'h00_00_ff;
            endcase
        end
        else begin  // JET
            case ( in_data )
            8'h00:  out_data = 24'h80_00_00;
            8'h01:  out_data = 24'h84_00_00;
            8'h02:  out_data = 24'h88_00_00;
            8'h03:  out_data = 24'h8c_00_00;
            8'h04:  out_data = 24'h90_00_00;
            8'h05:  out_data = 24'h94_00_00;
            8'h06:  out_data = 24'h98_00_00;
            8'h07:  out_data = 24'h9c_00_00;
            8'h08:  out_data = 24'ha0_00_00;
            8'h09:  out_data = 24'ha4_00_00;
            8'h0a:  out_data = 24'ha8_00_00;
            8'h0b:  out_data = 24'hac_00_00;
            8'h0c:  out_data = 24'hb0_00_00;
            8'h0d:  out_data = 24'hb4_00_00;
            8'h0e:  out_data = 24'hb8_00_00;
            8'h0f:  out_data = 24'hbc_00_00;
            8'h10:  out_data = 24'hc0_00_00;
            8'h11:  out_data = 24'hc4_00_00;
            8'h12:  out_data = 24'hc8_00_00;
            8'h13:  out_data = 24'hcc_00_00;
            8'h14:  out_data = 24'hd0_00_00;
            8'h15:  out_data = 24'hd4_00_00;
            8'h16:  out_data = 24'hd8_00_00;
            8'h17:  out_data = 24'hdc_00_00;
            8'h18:  out_data = 24'he0_00_00;
            8'h19:  out_data = 24'he4_00_00;
            8'h1a:  out_data = 24'he8_00_00;
            8'h1b:  out_data = 24'hec_00_00;
            8'h1c:  out_data = 24'hf0_00_00;
            8'h1d:  out_data = 24'hf4_00_00;
            8'h1e:  out_data = 24'hf8_00_00;
            8'h1f:  out_data = 24'hfc_00_00;
            8'h20:  out_data = 24'hff_00_00;
            8'h21:  out_data = 24'hff_04_00;
            8'h22:  out_data = 24'hff_08_00;
            8'h23:  out_data = 24'hff_0c_00;
            8'h24:  out_data = 24'hff_10_00;
            8'h25:  out_data = 24'hff_14_00;
            8'h26:  out_data = 24'hff_18_00;
            8'h27:  out_data = 24'hff_1c_00;
            8'h28:  out_data = 24'hff_20_00;
            8'h29:  out_data = 24'hff_24_00;
            8'h2a:  out_data = 24'hff_28_00;
            8'h2b:  out_data = 24'hff_2c_00;
            8'h2c:  out_data = 24'hff_30_00;
            8'h2d:  out_data = 24'hff_34_00;
            8'h2e:  out_data = 24'hff_38_00;
            8'h2f:  out_data = 24'hff_3c_00;
            8'h30:  out_data = 24'hff_40_00;
            8'h31:  out_data = 24'hff_44_00;
            8'h32:  out_data = 24'hff_48_00;
            8'h33:  out_data = 24'hff_4c_00;
            8'h34:  out_data = 24'hff_50_00;
            8'h35:  out_data = 24'hff_54_00;
            8'h36:  out_data = 24'hff_58_00;
            8'h37:  out_data = 24'hff_5c_00;
            8'h38:  out_data = 24'hff_60_00;
            8'h39:  out_data = 24'hff_64_00;
            8'h3a:  out_data = 24'hff_68_00;
            8'h3b:  out_data = 24'hff_6c_00;
            8'h3c:  out_data = 24'hff_70_00;
            8'h3d:  out_data = 24'hff_74_00;
            8'h3e:  out_data = 24'hff_78_00;
            8'h3f:  out_data = 24'hff_7c_00;
            8'h40:  out_data = 24'hff_80_00;
            8'h41:  out_data = 24'hff_84_00;
            8'h42:  out_data = 24'hff_88_00;
            8'h43:  out_data = 24'hff_8c_00;
            8'h44:  out_data = 24'hff_90_00;
            8'h45:  out_data = 24'hff_94_00;
            8'h46:  out_data = 24'hff_98_00;
            8'h47:  out_data = 24'hff_9c_00;
            8'h48:  out_data = 24'hff_a0_00;
            8'h49:  out_data = 24'hff_a4_00;
            8'h4a:  out_data = 24'hff_a8_00;
            8'h4b:  out_data = 24'hff_ac_00;
            8'h4c:  out_data = 24'hff_b0_00;
            8'h4d:  out_data = 24'hff_b4_00;
            8'h4e:  out_data = 24'hff_b8_00;
            8'h4f:  out_data = 24'hff_bc_00;
            8'h50:  out_data = 24'hff_c0_00;
            8'h51:  out_data = 24'hff_c4_00;
            8'h52:  out_data = 24'hff_c8_00;
            8'h53:  out_data = 24'hff_cc_00;
            8'h54:  out_data = 24'hff_d0_00;
            8'h55:  out_data = 24'hff_d4_00;
            8'h56:  out_data = 24'hff_d8_00;
            8'h57:  out_data = 24'hff_dc_00;
            8'h58:  out_data = 24'hff_e0_00;
            8'h59:  out_data = 24'hff_e4_00;
            8'h5a:  out_data = 24'hff_e8_00;
            8'h5b:  out_data = 24'hff_ec_00;
            8'h5c:  out_data = 24'hff_f0_00;
            8'h5d:  out_data = 24'hff_f4_00;
            8'h5e:  out_data = 24'hff_f8_00;
            8'h5f:  out_data = 24'hff_fc_00;
            8'h60:  out_data = 24'hfe_ff_02;
            8'h61:  out_data = 24'hfa_ff_06;
            8'h62:  out_data = 24'hf6_ff_0a;
            8'h63:  out_data = 24'hf2_ff_0e;
            8'h64:  out_data = 24'hee_ff_12;
            8'h65:  out_data = 24'hea_ff_16;
            8'h66:  out_data = 24'he6_ff_1a;
            8'h67:  out_data = 24'he2_ff_1e;
            8'h68:  out_data = 24'hde_ff_22;
            8'h69:  out_data = 24'hda_ff_26;
            8'h6a:  out_data = 24'hd6_ff_2a;
            8'h6b:  out_data = 24'hd2_ff_2e;
            8'h6c:  out_data = 24'hce_ff_32;
            8'h6d:  out_data = 24'hca_ff_36;
            8'h6e:  out_data = 24'hc6_ff_3a;
            8'h6f:  out_data = 24'hc2_ff_3e;
            8'h70:  out_data = 24'hbe_ff_42;
            8'h71:  out_data = 24'hba_ff_46;
            8'h72:  out_data = 24'hb6_ff_4a;
            8'h73:  out_data = 24'hb2_ff_4e;
            8'h74:  out_data = 24'hae_ff_52;
            8'h75:  out_data = 24'haa_ff_56;
            8'h76:  out_data = 24'ha6_ff_5a;
            8'h77:  out_data = 24'ha2_ff_5e;
            8'h78:  out_data = 24'h9e_ff_62;
            8'h79:  out_data = 24'h9a_ff_66;
            8'h7a:  out_data = 24'h96_ff_6a;
            8'h7b:  out_data = 24'h92_ff_6e;
            8'h7c:  out_data = 24'h8e_ff_72;
            8'h7d:  out_data = 24'h8a_ff_76;
            8'h7e:  out_data = 24'h86_ff_7a;
            8'h7f:  out_data = 24'h82_ff_7e;
            8'h80:  out_data = 24'h7e_ff_82;
            8'h81:  out_data = 24'h7a_ff_86;
            8'h82:  out_data = 24'h76_ff_8a;
            8'h83:  out_data = 24'h72_ff_8e;
            8'h84:  out_data = 24'h6e_ff_92;
            8'h85:  out_data = 24'h6a_ff_96;
            8'h86:  out_data = 24'h66_ff_9a;
            8'h87:  out_data = 24'h62_ff_9e;
            8'h88:  out_data = 24'h5e_ff_a2;
            8'h89:  out_data = 24'h5a_ff_a6;
            8'h8a:  out_data = 24'h56_ff_aa;
            8'h8b:  out_data = 24'h52_ff_ae;
            8'h8c:  out_data = 24'h4e_ff_b2;
            8'h8d:  out_data = 24'h4a_ff_b6;
            8'h8e:  out_data = 24'h46_ff_ba;
            8'h8f:  out_data = 24'h42_ff_be;
            8'h90:  out_data = 24'h3e_ff_c2;
            8'h91:  out_data = 24'h3a_ff_c6;
            8'h92:  out_data = 24'h36_ff_ca;
            8'h93:  out_data = 24'h32_ff_ce;
            8'h94:  out_data = 24'h2e_ff_d2;
            8'h95:  out_data = 24'h2a_ff_d6;
            8'h96:  out_data = 24'h26_ff_da;
            8'h97:  out_data = 24'h22_ff_de;
            8'h98:  out_data = 24'h1e_ff_e2;
            8'h99:  out_data = 24'h1a_ff_e6;
            8'h9a:  out_data = 24'h16_ff_ea;
            8'h9b:  out_data = 24'h12_ff_ee;
            8'h9c:  out_data = 24'h0e_ff_f2;
            8'h9d:  out_data = 24'h0a_ff_f6;
            8'h9e:  out_data = 24'h06_ff_fa;
            8'h9f:  out_data = 24'h01_ff_fe;
            8'ha0:  out_data = 24'h00_fc_ff;
            8'ha1:  out_data = 24'h00_f8_ff;
            8'ha2:  out_data = 24'h00_f4_ff;
            8'ha3:  out_data = 24'h00_f0_ff;
            8'ha4:  out_data = 24'h00_ec_ff;
            8'ha5:  out_data = 24'h00_e8_ff;
            8'ha6:  out_data = 24'h00_e4_ff;
            8'ha7:  out_data = 24'h00_e0_ff;
            8'ha8:  out_data = 24'h00_dc_ff;
            8'ha9:  out_data = 24'h00_d8_ff;
            8'haa:  out_data = 24'h00_d4_ff;
            8'hab:  out_data = 24'h00_d0_ff;
            8'hac:  out_data = 24'h00_cc_ff;
            8'had:  out_data = 24'h00_c8_ff;
            8'hae:  out_data = 24'h00_c4_ff;
            8'haf:  out_data = 24'h00_c0_ff;
            8'hb0:  out_data = 24'h00_bc_ff;
            8'hb1:  out_data = 24'h00_b8_ff;
            8'hb2:  out_data = 24'h00_b4_ff;
            8'hb3:  out_data = 24'h00_b0_ff;
            8'hb4:  out_data = 24'h00_ac_ff;
            8'hb5:  out_data = 24'h00_a8_ff;
            8'hb6:  out_data = 24'h00_a4_ff;
            8'hb7:  out_data = 24'h00_a0_ff;
            8'hb8:  out_data = 24'h00_9c_ff;
            8'hb9:  out_data = 24'h00_98_ff;
            8'hba:  out_data = 24'h00_94_ff;
            8'hbb:  out_data = 24'h00_90_ff;
            8'hbc:  out_data = 24'h00_8c_ff;
            8'hbd:  out_data = 24'h00_88_ff;
            8'hbe:  out_data = 24'h00_84_ff;
            8'hbf:  out_data = 24'h00_80_ff;
            8'hc0:  out_data = 24'h00_7c_ff;
            8'hc1:  out_data = 24'h00_78_ff;
            8'hc2:  out_data = 24'h00_74_ff;
            8'hc3:  out_data = 24'h00_70_ff;
            8'hc4:  out_data = 24'h00_6c_ff;
            8'hc5:  out_data = 24'h00_68_ff;
            8'hc6:  out_data = 24'h00_64_ff;
            8'hc7:  out_data = 24'h00_60_ff;
            8'hc8:  out_data = 24'h00_5c_ff;
            8'hc9:  out_data = 24'h00_58_ff;
            8'hca:  out_data = 24'h00_54_ff;
            8'hcb:  out_data = 24'h00_50_ff;
            8'hcc:  out_data = 24'h00_4c_ff;
            8'hcd:  out_data = 24'h00_48_ff;
            8'hce:  out_data = 24'h00_44_ff;
            8'hcf:  out_data = 24'h00_40_ff;
            8'hd0:  out_data = 24'h00_3c_ff;
            8'hd1:  out_data = 24'h00_38_ff;
            8'hd2:  out_data = 24'h00_34_ff;
            8'hd3:  out_data = 24'h00_30_ff;
            8'hd4:  out_data = 24'h00_2c_ff;
            8'hd5:  out_data = 24'h00_28_ff;
            8'hd6:  out_data = 24'h00_24_ff;
            8'hd7:  out_data = 24'h00_20_ff;
            8'hd8:  out_data = 24'h00_1c_ff;
            8'hd9:  out_data = 24'h00_18_ff;
            8'hda:  out_data = 24'h00_14_ff;
            8'hdb:  out_data = 24'h00_10_ff;
            8'hdc:  out_data = 24'h00_0c_ff;
            8'hdd:  out_data = 24'h00_08_ff;
            8'hde:  out_data = 24'h00_04_ff;
            8'hdf:  out_data = 24'h00_00_ff;
            8'he0:  out_data = 24'h00_00_fc;
            8'he1:  out_data = 24'h00_00_f8;
            8'he2:  out_data = 24'h00_00_f4;
            8'he3:  out_data = 24'h00_00_f0;
            8'he4:  out_data = 24'h00_00_ec;
            8'he5:  out_data = 24'h00_00_e8;
            8'he6:  out_data = 24'h00_00_e4;
            8'he7:  out_data = 24'h00_00_e0;
            8'he8:  out_data = 24'h00_00_dc;
            8'he9:  out_data = 24'h00_00_d8;
            8'hea:  out_data = 24'h00_00_d4;
            8'heb:  out_data = 24'h00_00_d0;
            8'hec:  out_data = 24'h00_00_cc;
            8'hed:  out_data = 24'h00_00_c8;
            8'hee:  out_data = 24'h00_00_c4;
            8'hef:  out_data = 24'h00_00_c0;
            8'hf0:  out_data = 24'h00_00_bc;
            8'hf1:  out_data = 24'h00_00_b8;
            8'hf2:  out_data = 24'h00_00_b4;
            8'hf3:  out_data = 24'h00_00_b0;
            8'hf4:  out_data = 24'h00_00_ac;
            8'hf5:  out_data = 24'h00_00_a8;
            8'hf6:  out_data = 24'h00_00_a4;
            8'hf7:  out_data = 24'h00_00_a0;
            8'hf8:  out_data = 24'h00_00_9c;
            8'hf9:  out_data = 24'h00_00_98;
            8'hfa:  out_data = 24'h00_00_94;
            8'hfb:  out_data = 24'h00_00_90;
            8'hfc:  out_data = 24'h00_00_8c;
            8'hfd:  out_data = 24'h00_00_88;
            8'hfe:  out_data = 24'h00_00_84;
            8'hff:  out_data = 24'h00_00_80;
            endcase
        end
    end
    
    
endmodule


`default_nettype wire


// end of file
