// ---------------------------------------------------------------------------
//  Jelly  -- the system on fpga system
//
//                                 Copyright (C) 2008-2016 by Ryuji Fuchikami
//                                 http://ryuz.my.coocan.jp/
//                                 https://github.com/ryuz/jelly.git
// ---------------------------------------------------------------------------



`timescale 1ns / 1ps
`default_nettype none



// multiplexer
module jelly_data_multiplexer
		#(
			parameter	NUM        = 5,
			parameter	DATA_WIDTH = 8,
			parameter	M_REGS     = 1
		)
		(
			input	wire							reset,
			input	wire							clk,
			input	wire							cke,
			
			input	wire							endian,
			
			input	wire	[NUM*DATA_WIDTH-1:0]	s_data,
			input	wire							s_valid,
			output	wire							s_ready,
			
			output	wire	[DATA_WIDTH-1:0]		m_data,
			output	wire							m_valid,
			input	wire							m_ready
		);
	
	localparam	SEL_WIDTH = NUM <=     2 ?  1 :
	                        NUM <=     4 ?  2 :
	                        NUM <=     8 ?  3 :
	                        NUM <=    16 ?  4 :
	                        NUM <=    32 ?  5 :
	                        NUM <=    64 ?  6 :
	                        NUM <=   128 ?  7 :
	                        NUM <=   256 ?  8 :
	                        NUM <=   512 ?  9 :
	                        NUM <=  1024 ? 10 :
	                        NUM <=  2048 ? 11 :
	                        NUM <=  4096 ? 12 :
	                        NUM <=  8192 ? 13 :
	                        NUM <= 16384 ? 14 :
	                        NUM <= 32768 ? 15 : 16;
	
	
	wire	[0:0]					stage_cke;
	wire	[0:0]					stage_valid;
	wire	[0:0]					next_valid;
	wire	[NUM*DATA_WIDTH-1:0]		src_data;
	wire							src_valid;
	wire	[DATA_WIDTH-1:0]	sink_data;
	
	jelly_pipeline_control
			#(
				.PIPELINE_STAGES	(1),
				.S_DATA_WIDTH		(NUM*DATA_WIDTH),
				.M_DATA_WIDTH		(DATA_WIDTH),
				.AUTO_VALID			(0),
				.MASTER_IN_REGS		(M_REGS),
				.MASTER_OUT_REGS	(M_REGS)
			)
		i_pipeline_control
			(
				.reset				(reset),
				.clk				(clk),
				.cke				(cke),
				
				.s_data				(s_data),
				.s_valid			(s_valid),
				.s_ready			(s_ready),
				
				.m_data				(m_data),
				.m_valid			(m_valid),
				.m_ready			(m_ready),
				
				.stage_cke			(stage_cke),
				.stage_valid		(stage_valid),
				.next_valid			(next_valid),
				.src_data			(src_data),
				.src_valid			(src_valid),
				.sink_data			(sink_data),
				.buffered			()
			);
	
	wire	[DATA_WIDTH-1:0]		sig_dout;
	
	reg		[SEL_WIDTH-1:0]			reg_sel;
	reg		[DATA_WIDTH-1:0]		reg_data;
	
	jelly_multiplexer
			#(
				.SEL_WIDTH		(SEL_WIDTH),
				.NUM			(NUM),
				.OUT_WIDTH		(DATA_WIDTH)
			)
		i_multiplexer
			(
				.endian			(endian),
				
				.sel			(reg_sel),
				.din			(src_data),
				.dout			(sig_dout)
			);
	
	always @(posedge clk) begin
		if ( reset ) begin
			reg_sel  <= {SEL_WIDTH{1'b0}};
			reg_data <= {(NUM*DATA_WIDTH){1'bx}};
		end
		else begin
			if ( stage_cke[0] ) begin
				if ( src_valid || reg_sel != {SEL_WIDTH{1'b0}} ) begin
					reg_sel  <= reg_sel + 1'b1;
					if ( reg_sel == (NUM-1) ) begin
						reg_sel  <= {SEL_WIDTH{1'b0}};
					end
					
					reg_data <= sig_dout;
				end
			end
		end
	end
	
	assign next_valid[0] = (src_valid || (reg_sel != {SEL_WIDTH{1'b0}}));
	
	assign sink_data     = reg_data;
	
	
endmodule



`default_nettype wire


// end of file
