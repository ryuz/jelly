
`timescale 1ns / 1ps
`default_nettype none


module tb_axi4_dummy_slave();
    localparam RATE = 1000.0/100.0;
    
    initial begin
        $dumpfile("tb_axi4_dummy_slave.vcd");
        $dumpvars(0, tb_axi4_dummy_slave);
        
        #100000;
            $finish;
    end
    
    reg     aclk = 1'b1;
    always #(RATE/2.0)      aclk = ~aclk;
    
    reg     aresetn = 1'b0;
    initial #(RATE*100) aresetn = 1'b1;
    
    parameter   RAND_BUSY = 0;
    
    parameter   BYTE_WIDTH       = 8;
    parameter   AXI4_ID_WIDTH    = 6;
    parameter   AXI4_ADDR_WIDTH  = 32;
    parameter   AXI4_DATA_SIZE   = 4;
    parameter   AXI4_DATA_WIDTH  = (BYTE_WIDTH << AXI4_DATA_SIZE);
    parameter   AXI4_STRB_WIDTH  = AXI4_DATA_WIDTH / BYTE_WIDTH;
    parameter   AXI4_LEN_WIDTH   = 2; //8;
    parameter   AXI4_QOS_WIDTH   = 4;
    
    wire    [AXI4_ID_WIDTH-1:0]     axi4_awid;
    wire    [AXI4_ADDR_WIDTH-1:0]   axi4_awaddr;
    wire    [AXI4_LEN_WIDTH-1:0]    axi4_awlen;
    wire    [2:0]                   axi4_awsize;
    wire    [1:0]                   axi4_awburst;
    wire    [0:0]                   axi4_awlock;
    wire    [3:0]                   axi4_awcache;
    wire    [2:0]                   axi4_awprot;
    wire    [AXI4_QOS_WIDTH-1:0]    axi4_awqos;
    wire    [3:0]                   axi4_awregion;
    wire                            axi4_awvalid;
    wire                            axi4_awready;
    wire    [AXI4_DATA_WIDTH-1:0]   axi4_wdata;
    wire    [AXI4_STRB_WIDTH-1:0]   axi4_wstrb;
    wire                            axi4_wlast;
    wire                            axi4_wvalid;
    wire                            axi4_wready;
    wire    [AXI4_ID_WIDTH-1:0]     axi4_bid;
    wire    [1:0]                   axi4_bresp;
    wire                            axi4_bvalid;
    wire                            axi4_bready;
    
    
    jelly_axi4_master_write_model
            #(
                .BYTE_WIDTH         (BYTE_WIDTH),
                .AXI4_ID_WIDTH      (AXI4_ID_WIDTH),
                .AXI4_ADDR_WIDTH    (AXI4_ADDR_WIDTH),
                .AXI4_DATA_SIZE     (AXI4_DATA_SIZE),
                .AXI4_DATA_WIDTH    (AXI4_DATA_WIDTH),
                .AXI4_STRB_WIDTH    (AXI4_STRB_WIDTH),
                .AXI4_LEN_WIDTH     (AXI4_LEN_WIDTH),
                .AXI4_QOS_WIDTH     (AXI4_QOS_WIDTH),
                .RATE_AW            (RAND_BUSY ? 50 : 100),
                .RATE_W             (RAND_BUSY ? 50 : 100),
                .RATE_B             (RAND_BUSY ? 50 : 100),
                .SEED_RAND          (1),
                .SEED_LEN           (2)
            )
        i_axi4_master_write_model
            (
                .aresetn            (aresetn),
                .aclk               (aclk),
                
                .m_axi4_awid        (axi4_awid),
                .m_axi4_awaddr      (axi4_awaddr),
                .m_axi4_awlen       (axi4_awlen),
                .m_axi4_awsize      (axi4_awsize),
                .m_axi4_awburst     (axi4_awburst),
                .m_axi4_awlock      (axi4_awlock),
                .m_axi4_awcache     (axi4_awcache),
                .m_axi4_awprot      (axi4_awprot),
                .m_axi4_awqos       (axi4_awqos),
                .m_axi4_awregion    (axi4_awregion),
                .m_axi4_awvalid     (axi4_awvalid),
                .m_axi4_awready     (axi4_awready),
                .m_axi4_wdata       (axi4_wdata),
                .m_axi4_wstrb       (axi4_wstrb),
                .m_axi4_wlast       (axi4_wlast),
                .m_axi4_wvalid      (axi4_wvalid),
                .m_axi4_wready      (axi4_wready),
                .m_axi4_bid         (axi4_bid),
                .m_axi4_bresp       (axi4_bresp),
                .m_axi4_bvalid      (axi4_bvalid),
                .m_axi4_bready      (axi4_bready)
            );
    
    
    wire    [AXI4_ID_WIDTH-1:0]     axi4_arid;
    wire    [AXI4_ADDR_WIDTH-1:0]   axi4_araddr;
    wire    [AXI4_LEN_WIDTH-1:0]    axi4_arlen;
    wire    [2:0]                   axi4_arsize;
    wire    [1:0]                   axi4_arburst;
    wire    [0:0]                   axi4_arlock;
    wire    [3:0]                   axi4_arcache;
    wire    [2:0]                   axi4_arprot;
    wire    [AXI4_QOS_WIDTH-1:0]    axi4_arqos;
    wire    [3:0]                   axi4_arregion;
    wire                            axi4_arvalid;
    wire                            axi4_arready;
    wire    [AXI4_ID_WIDTH-1:0]     axi4_rid;
    wire    [AXI4_DATA_WIDTH-1:0]   axi4_rdata;
    wire    [1:0]                   axi4_rresp;
    wire                            axi4_rlast;
    wire                            axi4_rvalid;
    wire                            axi4_rready;
    
    jelly_axi4_master_read_model
            #(
                .BYTE_WIDTH         (BYTE_WIDTH),
                .AXI4_ID_WIDTH      (AXI4_ID_WIDTH),
                .AXI4_ADDR_WIDTH    (AXI4_ADDR_WIDTH),
                .AXI4_DATA_SIZE     (AXI4_DATA_SIZE),
                .AXI4_DATA_WIDTH    (AXI4_DATA_WIDTH),
                .AXI4_STRB_WIDTH    (AXI4_STRB_WIDTH),
                .AXI4_LEN_WIDTH     (AXI4_LEN_WIDTH),
                .AXI4_QOS_WIDTH     (AXI4_QOS_WIDTH),
                
                .RATE_AR            (RAND_BUSY ? 50 : 100),
                .RATE_R             (RAND_BUSY ? 50 : 100),
                .SEED_RAND          (999)
            )
        i_axi4_master_read_model
            (
                .aresetn            (aresetn),
                .aclk               (aclk),
                
                .m_axi4_arid        (axi4_arid),
                .m_axi4_araddr      (axi4_araddr),
                .m_axi4_arlen       (axi4_arlen),
                .m_axi4_arsize      (axi4_arsize),
                .m_axi4_arburst     (axi4_arburst),
                .m_axi4_arlock      (axi4_arlock),
                .m_axi4_arcache     (axi4_arcache),
                .m_axi4_arprot      (axi4_arprot),
                .m_axi4_arqos       (axi4_arqos),
                .m_axi4_arregion    (axi4_arregion),
                .m_axi4_arvalid     (axi4_arvalid),
                .m_axi4_arready     (axi4_arready),
                .m_axi4_rid         (axi4_rid),
                .m_axi4_rdata       (axi4_rdata),
                .m_axi4_rresp       (axi4_rresp),
                .m_axi4_rlast       (axi4_rlast),
                .m_axi4_rvalid      (axi4_rvalid),
                .m_axi4_rready      (axi4_rready)
            );
    
    jelly_axi4_dummy_slave
            #(
                .BYTE_WIDTH         (BYTE_WIDTH),
                .AXI4_ID_WIDTH      (AXI4_ID_WIDTH),
                .AXI4_ADDR_WIDTH    (AXI4_ADDR_WIDTH),
                .AXI4_DATA_SIZE     (AXI4_DATA_SIZE),
                .AXI4_DATA_WIDTH    (AXI4_DATA_WIDTH),
                .AXI4_STRB_WIDTH    (AXI4_STRB_WIDTH),
                .AXI4_LEN_WIDTH     (AXI4_LEN_WIDTH),
                .AXI4_QOS_WIDTH     (AXI4_QOS_WIDTH)
            )
        i_axi4_dummy_slave
            (
                .aresetn            (aresetn),
                .aclk               (aclk),
                
                .s_axi4_awid        (axi4_awid),
                .s_axi4_awaddr      (axi4_awaddr),
                .s_axi4_awlen       (axi4_awlen),
                .s_axi4_awsize      (axi4_awsize),
                .s_axi4_awburst     (axi4_awburst),
                .s_axi4_awlock      (axi4_awlock),
                .s_axi4_awcache     (axi4_awcache),
                .s_axi4_awprot      (axi4_awprot),
                .s_axi4_awqos       (axi4_awqos),
                .s_axi4_awregion    (axi4_awregion),
                .s_axi4_awvalid     (axi4_awvalid),
                .s_axi4_awready     (axi4_awready),
                .s_axi4_wdata       (axi4_wdata),
                .s_axi4_wstrb       (axi4_wstrb),
                .s_axi4_wlast       (axi4_wlast),
                .s_axi4_wvalid      (axi4_wvalid),
                .s_axi4_wready      (axi4_wready),
                .s_axi4_bid         (axi4_bid),
                .s_axi4_bresp       (axi4_bresp),
                .s_axi4_bvalid      (axi4_bvalid),
                .s_axi4_bready      (axi4_bready),
                .s_axi4_arid        (axi4_arid),
                .s_axi4_araddr      (axi4_araddr),
                .s_axi4_arlen       (axi4_arlen),
                .s_axi4_arsize      (axi4_arsize),
                .s_axi4_arburst     (axi4_arburst),
                .s_axi4_arlock      (axi4_arlock),
                .s_axi4_arcache     (axi4_arcache),
                .s_axi4_arprot      (axi4_arprot),
                .s_axi4_arqos       (axi4_arqos),
                .s_axi4_arregion    (axi4_arregion),
                .s_axi4_arvalid     (axi4_arvalid),
                .s_axi4_arready     (axi4_arready),
                .s_axi4_rid         (axi4_rid),
                .s_axi4_rdata       (axi4_rdata),
                .s_axi4_rresp       (axi4_rresp),
                .s_axi4_rlast       (axi4_rlast),
                .s_axi4_rvalid      (axi4_rvalid),
                .s_axi4_rready      (axi4_rready)
            );
    
    
endmodule


`default_nettype wire


// end of file
