`timescale 1ns / 1ps

module boot_rom
		(
			clk ,
			addr,
			data
		);
	
	input				clk;
	input	[11:0]		addr;
	output	[31:0]		data;
	
	reg		[31:0]		data;
	
	always @ ( posedge clk ) begin
		case ( addr )
		12'h0:		data <= 32'h00000000;
		12'h1:		data <= 32'h00000000;
		12'h2:		data <= 32'h3c1c0101;
		12'h3:		data <= 32'h279c8240;
		12'h4:		data <= 32'h3c080000;
		12'h5:		data <= 32'h25082e98;
		12'h6:		data <= 32'h8d1d0000;
		12'h7:		data <= 32'h3c080100;
		12'h8:		data <= 32'h25080244;
		12'h9:		data <= 32'h3c090100;
		12'ha:		data <= 32'h252928ec;
		12'hb:		data <= 32'h11090005;
		12'hc:		data <= 32'h00000000;
		12'hd:		data <= 32'had000000;
		12'he:		data <= 32'h21080004;
		12'hf:		data <= 32'h1509fffd;
		12'h10:		data <= 32'h00000000;
		12'h11:		data <= 32'h3c080100;
		12'h12:		data <= 32'h25080000;
		12'h13:		data <= 32'h3c090100;
		12'h14:		data <= 32'h25290244;
		12'h15:		data <= 32'h3c0a0000;
		12'h16:		data <= 32'h254a2eb8;
		12'h17:		data <= 32'h11090007;
		12'h18:		data <= 32'h00000000;
		12'h19:		data <= 32'h8d4b0000;
		12'h1a:		data <= 32'h214a0004;
		12'h1b:		data <= 32'had0b0000;
		12'h1c:		data <= 32'h21080004;
		12'h1d:		data <= 32'h1509fffb;
		12'h1e:		data <= 32'h00000000;
		12'h1f:		data <= 32'h3c080000;
		12'h20:		data <= 32'h25080190;
		12'h21:		data <= 32'h0100f809;
		12'h22:		data <= 32'h00000000;
		12'h23:		data <= 32'h08000000;
		12'h24:		data <= 32'h00000000;
		12'h25:		data <= 32'h00000000;
		12'h26:		data <= 32'h00000000;
		12'h27:		data <= 32'h00000000;
		12'h28:		data <= 32'h00000000;
		12'h29:		data <= 32'h00000000;
		12'h2a:		data <= 32'h00000000;
		12'h2b:		data <= 32'h00000000;
		12'h2c:		data <= 32'h00000000;
		12'h2d:		data <= 32'h00000000;
		12'h2e:		data <= 32'h00000000;
		12'h2f:		data <= 32'h00000000;
		12'h30:		data <= 32'h00000000;
		12'h31:		data <= 32'h00000000;
		12'h32:		data <= 32'h00000000;
		12'h33:		data <= 32'h00000000;
		12'h34:		data <= 32'h00000000;
		12'h35:		data <= 32'h00000000;
		12'h36:		data <= 32'h00000000;
		12'h37:		data <= 32'h00000000;
		12'h38:		data <= 32'h00000000;
		12'h39:		data <= 32'h00000000;
		12'h3a:		data <= 32'h00000000;
		12'h3b:		data <= 32'h00000000;
		12'h3c:		data <= 32'h00000000;
		12'h3d:		data <= 32'h00000000;
		12'h3e:		data <= 32'h00000000;
		12'h3f:		data <= 32'h00000000;
		12'h40:		data <= 32'h00000000;
		12'h41:		data <= 32'h00000000;
		12'h42:		data <= 32'h00000000;
		12'h43:		data <= 32'h00000000;
		12'h44:		data <= 32'h00000000;
		12'h45:		data <= 32'h00000000;
		12'h46:		data <= 32'h00000000;
		12'h47:		data <= 32'h00000000;
		12'h48:		data <= 32'h00000000;
		12'h49:		data <= 32'h00000000;
		12'h4a:		data <= 32'h00000000;
		12'h4b:		data <= 32'h00000000;
		12'h4c:		data <= 32'h00000000;
		12'h4d:		data <= 32'h00000000;
		12'h4e:		data <= 32'h00000000;
		12'h4f:		data <= 32'h00000000;
		12'h50:		data <= 32'h00000000;
		12'h51:		data <= 32'h00000000;
		12'h52:		data <= 32'h00000000;
		12'h53:		data <= 32'h00000000;
		12'h54:		data <= 32'h00000000;
		12'h55:		data <= 32'h00000000;
		12'h56:		data <= 32'h00000000;
		12'h57:		data <= 32'h00000000;
		12'h58:		data <= 32'h00000000;
		12'h59:		data <= 32'h00000000;
		12'h5a:		data <= 32'h00000000;
		12'h5b:		data <= 32'h00000000;
		12'h5c:		data <= 32'h00000000;
		12'h5d:		data <= 32'h00000000;
		12'h5e:		data <= 32'h00000000;
		12'h5f:		data <= 32'h00000000;
		12'h60:		data <= 32'h3c1a0000;
		12'h61:		data <= 32'h275a1ef8;
		12'h62:		data <= 32'h03400008;
		12'h63:		data <= 32'h00000000;
		12'h64:		data <= 32'h27bdffe8;
		12'h65:		data <= 32'hafbf0010;
		12'h66:		data <= 32'h0c000259;
		12'h67:		data <= 32'h00000000;
		12'h68:		data <= 32'h8fbf0010;
		12'h69:		data <= 32'h00001021;
		12'h6a:		data <= 32'h03e00008;
		12'h6b:		data <= 32'h27bd0018;
		12'h6c:		data <= 32'h3c040100;
		12'h6d:		data <= 32'h3c060100;
		12'h6e:		data <= 32'h27bdffe8;
		12'h6f:		data <= 32'h248426b4;
		12'h70:		data <= 32'h24051000;
		12'h71:		data <= 32'hafbf0010;
		12'h72:		data <= 32'h0c000245;
		12'h73:		data <= 32'h24c61698;
		12'h74:		data <= 32'h3c050100;
		12'h75:		data <= 32'h3c020100;
		12'h76:		data <= 32'h3c030100;
		12'h77:		data <= 32'h24a52698;
		12'h78:		data <= 32'h244226dc;
		12'h79:		data <= 32'h24631088;
		12'h7a:		data <= 32'haca20038;
		12'h7b:		data <= 32'h24630200;
		12'h7c:		data <= 32'h3c020100;
		12'h7d:		data <= 32'h24040200;
		12'h7e:		data <= 32'hac4328e8;
		12'h7f:		data <= 32'haca40034;
		12'h80:		data <= 32'h8fbf0010;
		12'h81:		data <= 32'h00000000;
		12'h82:		data <= 32'h03e00008;
		12'h83:		data <= 32'h27bd0018;
		12'h84:		data <= 32'h27bdffe8;
		12'h85:		data <= 32'hafbf0010;
		12'h86:		data <= 32'h0c000201;
		12'h87:		data <= 32'h00002021;
		12'h88:		data <= 32'h8fbf0010;
		12'h89:		data <= 32'h00002021;
		12'h8a:		data <= 32'h08000096;
		12'h8b:		data <= 32'h27bd0018;
		12'h8c:		data <= 32'h27bdffe8;
		12'h8d:		data <= 32'hafbf0010;
		12'h8e:		data <= 32'h0c000197;
		12'h8f:		data <= 32'h00000000;
		12'h90:		data <= 32'h0c0001a3;
		12'h91:		data <= 32'h00402021;
		12'h92:		data <= 32'h8fbf0010;
		12'h93:		data <= 32'h24040001;
		12'h94:		data <= 32'h08000233;
		12'h95:		data <= 32'h27bd0018;
		12'h96:		data <= 32'h27bdffb8;
		12'h97:		data <= 32'hafbf0044;
		12'h98:		data <= 32'h0c000195;
		12'h99:		data <= 32'hafb00040;
		12'h9a:		data <= 32'h27a4001c;
		12'h9b:		data <= 32'h24030024;
		12'h9c:		data <= 32'h24020003;
		12'h9d:		data <= 32'hafa30024;
		12'h9e:		data <= 32'h24100001;
		12'h9f:		data <= 32'hafa20020;
		12'ha0:		data <= 32'hafa0001c;
		12'ha1:		data <= 32'h0c000590;
		12'ha2:		data <= 32'hafa00028;
		12'ha3:		data <= 32'h27a40010;
		12'ha4:		data <= 32'h3c030100;
		12'ha5:		data <= 32'hafb00014;
		12'ha6:		data <= 32'hac6228e0;
		12'ha7:		data <= 32'hafa00010;
		12'ha8:		data <= 32'h0c000414;
		12'ha9:		data <= 32'hafa00018;
		12'haa:		data <= 32'h3c030100;
		12'hab:		data <= 32'h24040001;
		12'hac:		data <= 32'h0c000298;
		12'had:		data <= 32'hac6228dc;
		12'hae:		data <= 32'h0c000298;
		12'haf:		data <= 32'h24040002;
		12'hb0:		data <= 32'h0c000298;
		12'hb1:		data <= 32'h24040003;
		12'hb2:		data <= 32'h0c000298;
		12'hb3:		data <= 32'h24040004;
		12'hb4:		data <= 32'h0c000298;
		12'hb5:		data <= 32'h24040005;
		12'hb6:		data <= 32'h0c000298;
		12'hb7:		data <= 32'h24040006;
		12'hb8:		data <= 32'h3c020000;
		12'hb9:		data <= 32'h27a4002c;
		12'hba:		data <= 32'h24420230;
		12'hbb:		data <= 32'hafb00034;
		12'hbc:		data <= 32'hafa20038;
		12'hbd:		data <= 32'hafa0002c;
		12'hbe:		data <= 32'h0c000706;
		12'hbf:		data <= 32'hafa00030;
		12'hc0:		data <= 32'h0c000221;
		12'hc1:		data <= 32'h24040001;
		12'hc2:		data <= 32'h8fbf0044;
		12'hc3:		data <= 32'h8fb00040;
		12'hc4:		data <= 32'h03e00008;
		12'hc5:		data <= 32'h27bd0048;
		12'hc6:		data <= 32'h27bdffe8;
		12'hc7:		data <= 32'h24040006;
		12'hc8:		data <= 32'hafbf0014;
		12'hc9:		data <= 32'h0c00039d;
		12'hca:		data <= 32'hafb00010;
		12'hcb:		data <= 32'h3c030100;
		12'hcc:		data <= 32'h8c700240;
		12'hcd:		data <= 32'h3c02015a;
		12'hce:		data <= 32'h34424e35;
		12'hcf:		data <= 32'h02020018;
		12'hd0:		data <= 32'h24040006;
		12'hd1:		data <= 32'h00008012;
		12'hd2:		data <= 32'h26100001;
		12'hd3:		data <= 32'h0c000343;
		12'hd4:		data <= 32'hac700240;
		12'hd5:		data <= 32'h3c031062;
		12'hd6:		data <= 32'h34634dd3;
		12'hd7:		data <= 32'h02030019;
		12'hd8:		data <= 32'h8fbf0014;
		12'hd9:		data <= 32'h00001810;
		12'hda:		data <= 32'h00031982;
		12'hdb:		data <= 32'h00032080;
		12'hdc:		data <= 32'h000311c0;
		12'hdd:		data <= 32'h00441023;
		12'hde:		data <= 32'h00431021;
		12'hdf:		data <= 32'h000210c0;
		12'he0:		data <= 32'h02028023;
		12'he1:		data <= 32'h26040064;
		12'he2:		data <= 32'h8fb00010;
		12'he3:		data <= 32'h080002ff;
		12'he4:		data <= 32'h27bd0018;
		12'he5:		data <= 32'h27bdffd8;
		12'he6:		data <= 32'hafb1001c;
		12'he7:		data <= 32'hafb00018;
		12'he8:		data <= 32'hafbf0020;
		12'he9:		data <= 32'h3c020100;
		12'hea:		data <= 32'h00808021;
		12'heb:		data <= 32'h8c4428e0;
		12'hec:		data <= 32'h00a08821;
		12'hed:		data <= 32'h0c000616;
		12'hee:		data <= 32'h27a50010;
		12'hef:		data <= 32'h8fa50010;
		12'hf0:		data <= 32'h24030020;
		12'hf1:		data <= 32'h2402003a;
		12'hf2:		data <= 32'h26100030;
		12'hf3:		data <= 32'ha0b00004;
		12'hf4:		data <= 32'ha0a20006;
		12'hf5:		data <= 32'ha0a30007;
		12'hf6:		data <= 32'ha0a30005;
		12'hf7:		data <= 32'h82220000;
		12'hf8:		data <= 32'h00000000;
		12'hf9:		data <= 32'h14400011;
		12'hfa:		data <= 32'h00a01821;
		12'hfb:		data <= 32'h24020004;
		12'hfc:		data <= 32'h24060005;
		12'hfd:		data <= 32'h00a21821;
		12'hfe:		data <= 32'h00a62021;
		12'hff:		data <= 32'h2402000a;
		12'h100:		data <= 32'ha0620004;
		12'h101:		data <= 32'ha0800004;
		12'h102:		data <= 32'h3c020100;
		12'h103:		data <= 32'h8c4428dc;
		12'h104:		data <= 32'h0c0004ae;
		12'h105:		data <= 32'h00000000;
		12'h106:		data <= 32'h8fbf0020;
		12'h107:		data <= 32'h8fb1001c;
		12'h108:		data <= 32'h8fb00018;
		12'h109:		data <= 32'h03e00008;
		12'h10a:		data <= 32'h27bd0028;
		12'h10b:		data <= 32'h00002021;
		12'h10c:		data <= 32'h24840001;
		12'h10d:		data <= 32'ha0620008;
		12'h10e:		data <= 32'h02241021;
		12'h10f:		data <= 32'h80420000;
		12'h110:		data <= 32'h00000000;
		12'h111:		data <= 32'h1440fffa;
		12'h112:		data <= 32'h24630001;
		12'h113:		data <= 32'h24820004;
		12'h114:		data <= 32'h24860005;
		12'h115:		data <= 32'h00a21821;
		12'h116:		data <= 32'h00a62021;
		12'h117:		data <= 32'h2402000a;
		12'h118:		data <= 32'ha0620004;
		12'h119:		data <= 32'ha0800004;
		12'h11a:		data <= 32'h3c020100;
		12'h11b:		data <= 32'h8c4428dc;
		12'h11c:		data <= 32'h0c0004ae;
		12'h11d:		data <= 32'h00000000;
		12'h11e:		data <= 32'h8fbf0020;
		12'h11f:		data <= 32'h8fb1001c;
		12'h120:		data <= 32'h8fb00018;
		12'h121:		data <= 32'h03e00008;
		12'h122:		data <= 32'h27bd0028;
		12'h123:		data <= 32'h27bdffc8;
		12'h124:		data <= 32'hafb7002c;
		12'h125:		data <= 32'hafb60028;
		12'h126:		data <= 32'hafb50024;
		12'h127:		data <= 32'hafb40020;
		12'h128:		data <= 32'hafb3001c;
		12'h129:		data <= 32'hafb20018;
		12'h12a:		data <= 32'hafb10014;
		12'h12b:		data <= 32'hafb00010;
		12'h12c:		data <= 32'hafbf0030;
		12'h12d:		data <= 32'h0080a021;
		12'h12e:		data <= 32'h3c170000;
		12'h12f:		data <= 32'h28910002;
		12'h130:		data <= 32'h2492ffff;
		12'h131:		data <= 32'h28900005;
		12'h132:		data <= 32'h24930001;
		12'h133:		data <= 32'h3c150000;
		12'h134:		data <= 32'h3c160000;
		12'h135:		data <= 32'h02802021;
		12'h136:		data <= 32'h0c0000e5;
		12'h137:		data <= 32'h26e52e9c;
		12'h138:		data <= 32'h0c0000c6;
		12'h139:		data <= 32'h00000000;
		12'h13a:		data <= 32'h0800015f;
		12'h13b:		data <= 32'h00000000;
		12'h13c:		data <= 32'h0c00039f;
		12'h13d:		data <= 32'h24040001;
		12'h13e:		data <= 32'h1040002b;
		12'h13f:		data <= 32'h02802021;
		12'h140:		data <= 32'h16200002;
		12'h141:		data <= 32'h24040005;
		12'h142:		data <= 32'h02402021;
		12'h143:		data <= 32'h0c000343;
		12'h144:		data <= 32'h00000000;
		12'h145:		data <= 32'h02802021;
		12'h146:		data <= 32'h0c0000e5;
		12'h147:		data <= 32'h26a52ea8;
		12'h148:		data <= 32'h0c0000c6;
		12'h149:		data <= 32'h00000000;
		12'h14a:		data <= 32'h1600002e;
		12'h14b:		data <= 32'h00000000;
		12'h14c:		data <= 32'h0c00039d;
		12'h14d:		data <= 32'h24040001;
		12'h14e:		data <= 32'h16200002;
		12'h14f:		data <= 32'h24040005;
		12'h150:		data <= 32'h02402021;
		12'h151:		data <= 32'h0c00039f;
		12'h152:		data <= 32'h00000000;
		12'h153:		data <= 32'h10400016;
		12'h154:		data <= 32'h02802021;
		12'h155:		data <= 32'h16000002;
		12'h156:		data <= 32'h02602021;
		12'h157:		data <= 32'h24040001;
		12'h158:		data <= 32'h0c000343;
		12'h159:		data <= 32'h00000000;
		12'h15a:		data <= 32'h02802021;
		12'h15b:		data <= 32'h0c0000e5;
		12'h15c:		data <= 32'h26a52ea8;
		12'h15d:		data <= 32'h0c0000c6;
		12'h15e:		data <= 32'h00000000;
		12'h15f:		data <= 32'h16200002;
		12'h160:		data <= 32'h24040005;
		12'h161:		data <= 32'h02402021;
		12'h162:		data <= 32'h0c00039d;
		12'h163:		data <= 32'h00000000;
		12'h164:		data <= 32'h1200ffd7;
		12'h165:		data <= 32'h00000000;
		12'h166:		data <= 32'h0c00039f;
		12'h167:		data <= 32'h02602021;
		12'h168:		data <= 32'h1440ffd7;
		12'h169:		data <= 32'h02802021;
		12'h16a:		data <= 32'h0c0000e5;
		12'h16b:		data <= 32'h26c52eb0;
		12'h16c:		data <= 32'h0c0000c6;
		12'h16d:		data <= 32'h00000000;
		12'h16e:		data <= 32'h16200002;
		12'h16f:		data <= 32'h24040005;
		12'h170:		data <= 32'h02402021;
		12'h171:		data <= 32'h0c000343;
		12'h172:		data <= 32'h00000000;
		12'h173:		data <= 32'h1600000b;
		12'h174:		data <= 32'h00000000;
		12'h175:		data <= 32'h0c000343;
		12'h176:		data <= 32'h24040001;
		12'h177:		data <= 32'h08000136;
		12'h178:		data <= 32'h02802021;
		12'h179:		data <= 32'h0c00039d;
		12'h17a:		data <= 32'h02602021;
		12'h17b:		data <= 32'h1220ffd4;
		12'h17c:		data <= 32'h24040005;
		12'h17d:		data <= 32'h08000151;
		12'h17e:		data <= 32'h00000000;
		12'h17f:		data <= 32'h0c000343;
		12'h180:		data <= 32'h02602021;
		12'h181:		data <= 32'h08000136;
		12'h182:		data <= 32'h02802021;
		12'h183:		data <= 32'h27bdffd8;
		12'h184:		data <= 32'hafb1001c;
		12'h185:		data <= 32'hafb00018;
		12'h186:		data <= 32'hafbf0020;
		12'h187:		data <= 32'h3c110100;
		12'h188:		data <= 32'h3c100100;
		12'h189:		data <= 32'h8e2428dc;
		12'h18a:		data <= 32'h0c0004ed;
		12'h18b:		data <= 32'h27a50010;
		12'h18c:		data <= 32'h8fa40010;
		12'h18d:		data <= 32'h0c0001ad;
		12'h18e:		data <= 32'h24840004;
		12'h18f:		data <= 32'h8e0428e0;
		12'h190:		data <= 32'h8fa50010;
		12'h191:		data <= 32'h0c00067a;
		12'h192:		data <= 32'h00000000;
		12'h193:		data <= 32'h08000189;
		12'h194:		data <= 32'h00000000;
		12'h195:		data <= 32'h03e00008;
		12'h196:		data <= 32'h00000000;
		12'h197:		data <= 32'h3c04f200;
		12'h198:		data <= 32'h34830004;
		12'h199:		data <= 32'h8c620000;
		12'h19a:		data <= 32'h00000000;
		12'h19b:		data <= 32'h30420001;
		12'h19c:		data <= 32'h1040fffc;
		12'h19d:		data <= 32'h00000000;
		12'h19e:		data <= 32'h8c820000;
		12'h19f:		data <= 32'h00000000;
		12'h1a0:		data <= 32'h00021600;
		12'h1a1:		data <= 32'h03e00008;
		12'h1a2:		data <= 32'h00021603;
		12'h1a3:		data <= 32'h3c05f200;
		12'h1a4:		data <= 32'h34a30004;
		12'h1a5:		data <= 32'h8c620000;
		12'h1a6:		data <= 32'h00000000;
		12'h1a7:		data <= 32'h30420002;
		12'h1a8:		data <= 32'h1040fffc;
		12'h1a9:		data <= 32'h00000000;
		12'h1aa:		data <= 32'haca40000;
		12'h1ab:		data <= 32'h03e00008;
		12'h1ac:		data <= 32'h00000000;
		12'h1ad:		data <= 32'h27bdffe0;
		12'h1ae:		data <= 32'hafb00010;
		12'h1af:		data <= 32'hafbf0018;
		12'h1b0:		data <= 32'hafb10014;
		12'h1b1:		data <= 32'h80820000;
		12'h1b2:		data <= 32'h00000000;
		12'h1b3:		data <= 32'h10400014;
		12'h1b4:		data <= 32'h00808021;
		12'h1b5:		data <= 32'h080001be;
		12'h1b6:		data <= 32'h2411000a;
		12'h1b7:		data <= 32'h00402021;
		12'h1b8:		data <= 32'h0c0001a3;
		12'h1b9:		data <= 32'h26100001;
		12'h1ba:		data <= 32'h82020000;
		12'h1bb:		data <= 32'h00000000;
		12'h1bc:		data <= 32'h1040000b;
		12'h1bd:		data <= 32'h00000000;
		12'h1be:		data <= 32'h1451fff8;
		12'h1bf:		data <= 32'h2404000d;
		12'h1c0:		data <= 32'h0c0001a3;
		12'h1c1:		data <= 32'h26100001;
		12'h1c2:		data <= 32'h0c0001a3;
		12'h1c3:		data <= 32'h2404000a;
		12'h1c4:		data <= 32'h82020000;
		12'h1c5:		data <= 32'h00000000;
		12'h1c6:		data <= 32'h1440fff7;
		12'h1c7:		data <= 32'h00000000;
		12'h1c8:		data <= 32'h8fbf0018;
		12'h1c9:		data <= 32'h8fb10014;
		12'h1ca:		data <= 32'h8fb00010;
		12'h1cb:		data <= 32'h03e00008;
		12'h1cc:		data <= 32'h27bd0020;
		12'h1cd:		data <= 32'h24820030;
		12'h1ce:		data <= 32'h00021600;
		12'h1cf:		data <= 32'h24830057;
		12'h1d0:		data <= 32'h2884000a;
		12'h1d1:		data <= 32'h14800003;
		12'h1d2:		data <= 32'h00021603;
		12'h1d3:		data <= 32'h00031600;
		12'h1d4:		data <= 32'h00021603;
		12'h1d5:		data <= 32'h03e00008;
		12'h1d6:		data <= 32'h00000000;
		12'h1d7:		data <= 32'h27bdffe8;
		12'h1d8:		data <= 32'hafb00010;
		12'h1d9:		data <= 32'h00048600;
		12'h1da:		data <= 32'h00108603;
		12'h1db:		data <= 32'h00102103;
		12'h1dc:		data <= 32'hafbf0014;
		12'h1dd:		data <= 32'h0c0001cd;
		12'h1de:		data <= 32'h3084000f;
		12'h1df:		data <= 32'h0c0001a3;
		12'h1e0:		data <= 32'h00402021;
		12'h1e1:		data <= 32'h0c0001cd;
		12'h1e2:		data <= 32'h3204000f;
		12'h1e3:		data <= 32'h00402021;
		12'h1e4:		data <= 32'h8fbf0014;
		12'h1e5:		data <= 32'h8fb00010;
		12'h1e6:		data <= 32'h080001a3;
		12'h1e7:		data <= 32'h27bd0018;
		12'h1e8:		data <= 32'h27bdffe8;
		12'h1e9:		data <= 32'hafb00010;
		12'h1ea:		data <= 32'h3090ffff;
		12'h1eb:		data <= 32'h00102202;
		12'h1ec:		data <= 32'h00042600;
		12'h1ed:		data <= 32'hafbf0014;
		12'h1ee:		data <= 32'h0c0001d7;
		12'h1ef:		data <= 32'h00042603;
		12'h1f0:		data <= 32'h00102600;
		12'h1f1:		data <= 32'h8fbf0014;
		12'h1f2:		data <= 32'h8fb00010;
		12'h1f3:		data <= 32'h00042603;
		12'h1f4:		data <= 32'h080001d7;
		12'h1f5:		data <= 32'h27bd0018;
		12'h1f6:		data <= 32'h27bdffe8;
		12'h1f7:		data <= 32'hafb00010;
		12'h1f8:		data <= 32'h00808021;
		12'h1f9:		data <= 32'hafbf0014;
		12'h1fa:		data <= 32'h0c0001e8;
		12'h1fb:		data <= 32'h00042402;
		12'h1fc:		data <= 32'h3204ffff;
		12'h1fd:		data <= 32'h8fbf0014;
		12'h1fe:		data <= 32'h8fb00010;
		12'h1ff:		data <= 32'h080001e8;
		12'h200:		data <= 32'h27bd0018;
		12'h201:		data <= 32'h27bdffd8;
		12'h202:		data <= 32'h3c020000;
		12'h203:		data <= 32'h27a40010;
		12'h204:		data <= 32'h24420868;
		12'h205:		data <= 32'hafbf0020;
		12'h206:		data <= 32'hafa2001c;
		12'h207:		data <= 32'hafa00010;
		12'h208:		data <= 32'hafa00014;
		12'h209:		data <= 32'h0c000706;
		12'h20a:		data <= 32'hafa00018;
		12'h20b:		data <= 32'h3c05f100;
		12'h20c:		data <= 32'h34a60004;
		12'h20d:		data <= 32'h3402c34f;
		12'h20e:		data <= 32'hacc20000;
		12'h20f:		data <= 32'h24030002;
		12'h210:		data <= 32'h24020001;
		12'h211:		data <= 32'haca30000;
		12'h212:		data <= 32'h00002021;
		12'h213:		data <= 32'haca20000;
		12'h214:		data <= 32'h0c000221;
		12'h215:		data <= 32'h00000000;
		12'h216:		data <= 32'h8fbf0020;
		12'h217:		data <= 32'h00000000;
		12'h218:		data <= 32'h03e00008;
		12'h219:		data <= 32'h27bd0028;
		12'h21a:		data <= 32'h27bdffe8;
		12'h21b:		data <= 32'hafbf0010;
		12'h21c:		data <= 32'h0c000233;
		12'h21d:		data <= 32'h00002021;
		12'h21e:		data <= 32'h8fbf0010;
		12'h21f:		data <= 32'h080006e7;
		12'h220:		data <= 32'h27bd0018;
		12'h221:		data <= 32'h3c03f000;
		12'h222:		data <= 32'h34620010;
		12'h223:		data <= 32'h04810004;
		12'h224:		data <= 32'h00802821;
		12'h225:		data <= 32'h2405ffef;
		12'h226:		data <= 32'h03e00008;
		12'h227:		data <= 32'h00a01021;
		12'h228:		data <= 32'h8c420000;
		12'h229:		data <= 32'h00042100;
		12'h22a:		data <= 32'h34630020;
		12'h22b:		data <= 32'h0045102b;
		12'h22c:		data <= 32'h00831821;
		12'h22d:		data <= 32'h1440fff7;
		12'h22e:		data <= 32'h00002821;
		12'h22f:		data <= 32'h24020001;
		12'h230:		data <= 32'hac620000;
		12'h231:		data <= 32'h03e00008;
		12'h232:		data <= 32'h00a01021;
		12'h233:		data <= 32'h3c03f000;
		12'h234:		data <= 32'h34620010;
		12'h235:		data <= 32'h04810004;
		12'h236:		data <= 32'h00802821;
		12'h237:		data <= 32'h2405ffef;
		12'h238:		data <= 32'h03e00008;
		12'h239:		data <= 32'h00a01021;
		12'h23a:		data <= 32'h8c420000;
		12'h23b:		data <= 32'h00042100;
		12'h23c:		data <= 32'h34630024;
		12'h23d:		data <= 32'h0045102b;
		12'h23e:		data <= 32'h00831821;
		12'h23f:		data <= 32'h1440fff7;
		12'h240:		data <= 32'h00002821;
		12'h241:		data <= 32'h00a01021;
		12'h242:		data <= 32'hac600000;
		12'h243:		data <= 32'h03e00008;
		12'h244:		data <= 32'h00000000;
		12'h245:		data <= 32'h2402ffe0;
		12'h246:		data <= 32'h00a22824;
		12'h247:		data <= 32'h00c54021;
		12'h248:		data <= 32'h2ca2000d;
		12'h249:		data <= 32'h24a9ffc0;
		12'h24a:		data <= 32'h10400003;
		12'h24b:		data <= 32'h2507ffe0;
		12'h24c:		data <= 32'h03e00008;
		12'h24d:		data <= 32'hac800000;
		12'h24e:		data <= 32'h3402abcd;
		12'h24f:		data <= 32'h24031234;
		12'h250:		data <= 32'hac850004;
		12'h251:		data <= 32'hac860000;
		12'h252:		data <= 32'hacc20008;
		12'h253:		data <= 32'hacc90004;
		12'h254:		data <= 32'hacc00000;
		12'h255:		data <= 32'hace30008;
		12'h256:		data <= 32'hace00004;
		12'h257:		data <= 32'h03e00008;
		12'h258:		data <= 32'had00ffe0;
		12'h259:		data <= 32'h27bdffd8;
		12'h25a:		data <= 32'hafb00018;
		12'h25b:		data <= 32'h3c100100;
		12'h25c:		data <= 32'h26102698;
		12'h25d:		data <= 32'hafbf0020;
		12'h25e:		data <= 32'h0c000786;
		12'h25f:		data <= 32'hafb1001c;
		12'h260:		data <= 32'h8e020024;
		12'h261:		data <= 32'h3c110100;
		12'h262:		data <= 32'h34420005;
		12'h263:		data <= 32'h0c0007fb;
		12'h264:		data <= 32'hae020024;
		12'h265:		data <= 32'h0c00006c;
		12'h266:		data <= 32'h00000000;
		12'h267:		data <= 32'h8e020038;
		12'h268:		data <= 32'h8e050034;
		12'h269:		data <= 32'h3c060000;
		12'h26a:		data <= 32'h00452821;
		12'h26b:		data <= 32'h24c60a0c;
		12'h26c:		data <= 32'h262426c8;
		12'h26d:		data <= 32'h00003821;
		12'h26e:		data <= 32'h0c000797;
		12'h26f:		data <= 32'hafa00010;
		12'h270:		data <= 32'h8e020024;
		12'h271:		data <= 32'h00000000;
		12'h272:		data <= 32'h30420009;
		12'h273:		data <= 32'h14400003;
		12'h274:		data <= 32'h00000000;
		12'h275:		data <= 32'h0c00078e;
		12'h276:		data <= 32'h00000000;
		12'h277:		data <= 32'h0c000084;
		12'h278:		data <= 32'h00000000;
		12'h279:		data <= 32'h0c000786;
		12'h27a:		data <= 32'h00000000;
		12'h27b:		data <= 32'h0c0007b0;
		12'h27c:		data <= 32'h262426c8;
		12'h27d:		data <= 32'h8fbf0020;
		12'h27e:		data <= 32'h8fb1001c;
		12'h27f:		data <= 32'h8fb00018;
		12'h280:		data <= 32'h00001021;
		12'h281:		data <= 32'h03e00008;
		12'h282:		data <= 32'h27bd0028;
		12'h283:		data <= 32'h27bdffe8;
		12'h284:		data <= 32'hafb00010;
		12'h285:		data <= 32'h3c100100;
		12'h286:		data <= 32'hafbf0014;
		12'h287:		data <= 32'h26102698;
		12'h288:		data <= 32'h8e020024;
		12'h289:		data <= 32'h2403fff0;
		12'h28a:		data <= 32'h00431024;
		12'h28b:		data <= 32'h0c00082b;
		12'h28c:		data <= 32'hae020024;
		12'h28d:		data <= 32'h8e020024;
		12'h28e:		data <= 32'h00000000;
		12'h28f:		data <= 32'h30420009;
		12'h290:		data <= 32'h14400003;
		12'h291:		data <= 32'h00000000;
		12'h292:		data <= 32'h0c00078e;
		12'h293:		data <= 32'h00000000;
		12'h294:		data <= 32'h8fbf0014;
		12'h295:		data <= 32'h8fb00010;
		12'h296:		data <= 32'h08000823;
		12'h297:		data <= 32'h27bd0018;
		12'h298:		data <= 32'h27bdffd8;
		12'h299:		data <= 32'hafb00018;
		12'h29a:		data <= 32'hafbf0020;
		12'h29b:		data <= 32'hafb1001c;
		12'h29c:		data <= 32'h1480000d;
		12'h29d:		data <= 32'h00808021;
		12'h29e:		data <= 32'h3c110100;
		12'h29f:		data <= 32'h26232698;
		12'h2a0:		data <= 32'h8c620024;
		12'h2a1:		data <= 32'h00000000;
		12'h2a2:		data <= 32'h30420004;
		12'h2a3:		data <= 32'h1040001a;
		12'h2a4:		data <= 32'h2402ffee;
		12'h2a5:		data <= 32'h8fbf0020;
		12'h2a6:		data <= 32'h8fb1001c;
		12'h2a7:		data <= 32'h8fb00018;
		12'h2a8:		data <= 32'h03e00008;
		12'h2a9:		data <= 32'h27bd0028;
		12'h2aa:		data <= 32'h1880fffa;
		12'h2ab:		data <= 32'h2402ffee;
		12'h2ac:		data <= 32'h3c030000;
		12'h2ad:		data <= 32'h8c622e94;
		12'h2ae:		data <= 32'h00000000;
		12'h2af:		data <= 32'h0044102a;
		12'h2b0:		data <= 32'h1440fff4;
		12'h2b1:		data <= 32'h2402ffee;
		12'h2b2:		data <= 32'h0c000786;
		12'h2b3:		data <= 32'h00000000;
		12'h2b4:		data <= 32'h3c050100;
		12'h2b5:		data <= 32'h00101080;
		12'h2b6:		data <= 32'h24a30078;
		12'h2b7:		data <= 32'h00431021;
		12'h2b8:		data <= 32'h8c44fffc;
		12'h2b9:		data <= 32'h00000000;
		12'h2ba:		data <= 32'h10800038;
		12'h2bb:		data <= 32'h3c110100;
		12'h2bc:		data <= 32'h080002c3;
		12'h2bd:		data <= 32'h24a20078;
		12'h2be:		data <= 32'h8c70002c;
		12'h2bf:		data <= 32'h0c000786;
		12'h2c0:		data <= 32'h00000000;
		12'h2c1:		data <= 32'h3c050100;
		12'h2c2:		data <= 32'h24a20078;
		12'h2c3:		data <= 32'h00101880;
		12'h2c4:		data <= 32'h00621821;
		12'h2c5:		data <= 32'h8c64fffc;
		12'h2c6:		data <= 32'h00000000;
		12'h2c7:		data <= 32'h90820018;
		12'h2c8:		data <= 32'h00000000;
		12'h2c9:		data <= 32'h10400015;
		12'h2ca:		data <= 32'h24020002;
		12'h2cb:		data <= 32'h9082001d;
		12'h2cc:		data <= 32'h00000000;
		12'h2cd:		data <= 32'h24420001;
		12'h2ce:		data <= 32'ha082001d;
		12'h2cf:		data <= 32'h26232698;
		12'h2d0:		data <= 32'h8c620024;
		12'h2d1:		data <= 32'h00000000;
		12'h2d2:		data <= 32'h30420009;
		12'h2d3:		data <= 32'h10400007;
		12'h2d4:		data <= 32'h00000000;
		12'h2d5:		data <= 32'h00001021;
		12'h2d6:		data <= 32'h8fbf0020;
		12'h2d7:		data <= 32'h8fb1001c;
		12'h2d8:		data <= 32'h8fb00018;
		12'h2d9:		data <= 32'h03e00008;
		12'h2da:		data <= 32'h27bd0028;
		12'h2db:		data <= 32'h0c00078e;
		12'h2dc:		data <= 32'h00000000;
		12'h2dd:		data <= 32'h080002d6;
		12'h2de:		data <= 32'h00001021;
		12'h2df:		data <= 32'h9083003c;
		12'h2e0:		data <= 32'h8c850040;
		12'h2e1:		data <= 32'h8c870034;
		12'h2e2:		data <= 32'h8c880038;
		12'h2e3:		data <= 32'h3c060000;
		12'h2e4:		data <= 32'ha083001a;
		12'h2e5:		data <= 32'ha0820018;
		12'h2e6:		data <= 32'ha0830019;
		12'h2e7:		data <= 32'ha080001d;
		12'h2e8:		data <= 32'ha080001e;
		12'h2e9:		data <= 32'ha080001f;
		12'h2ea:		data <= 32'h24c62040;
		12'h2eb:		data <= 32'h0c000797;
		12'h2ec:		data <= 32'hafa80010;
		12'h2ed:		data <= 32'h0c000869;
		12'h2ee:		data <= 32'h02002021;
		12'h2ef:		data <= 32'h0c00082b;
		12'h2f0:		data <= 32'h00000000;
		12'h2f1:		data <= 32'h080002d0;
		12'h2f2:		data <= 32'h26232698;
		12'h2f3:		data <= 32'h3c030100;
		12'h2f4:		data <= 32'h8c6226bc;
		12'h2f5:		data <= 32'h00000000;
		12'h2f6:		data <= 32'h30420009;
		12'h2f7:		data <= 32'h10400003;
		12'h2f8:		data <= 32'h00000000;
		12'h2f9:		data <= 32'h080002a5;
		12'h2fa:		data <= 32'h2402ffd6;
		12'h2fb:		data <= 32'h0c00078e;
		12'h2fc:		data <= 32'h00000000;
		12'h2fd:		data <= 32'h080002a5;
		12'h2fe:		data <= 32'h2402ffd6;
		12'h2ff:		data <= 32'h27bdffd8;
		12'h300:		data <= 32'h3c020100;
		12'h301:		data <= 32'hafb3001c;
		12'h302:		data <= 32'hafb20018;
		12'h303:		data <= 32'hafbf0020;
		12'h304:		data <= 32'h24522698;
		12'h305:		data <= 32'hafb10014;
		12'h306:		data <= 32'hafb00010;
		12'h307:		data <= 32'h8e51002c;
		12'h308:		data <= 32'h0c000786;
		12'h309:		data <= 32'h00809821;
		12'h30a:		data <= 32'h3c020100;
		12'h30b:		data <= 32'h24420078;
		12'h30c:		data <= 32'h00111880;
		12'h30d:		data <= 32'h00621821;
		12'h30e:		data <= 32'h8e420024;
		12'h30f:		data <= 32'h02202021;
		12'h310:		data <= 32'h1440002c;
		12'h311:		data <= 32'h30450009;
		12'h312:		data <= 32'h8c70fffc;
		12'h313:		data <= 32'h0c000874;
		12'h314:		data <= 32'h00000000;
		12'h315:		data <= 32'h24020004;
		12'h316:		data <= 32'h24030001;
		12'h317:		data <= 32'h3c040100;
		12'h318:		data <= 32'ha2020018;
		12'h319:		data <= 32'ha203001b;
		12'h31a:		data <= 32'h248426a4;
		12'h31b:		data <= 32'h02202821;
		12'h31c:		data <= 32'h0c000980;
		12'h31d:		data <= 32'h02603021;
		12'h31e:		data <= 32'h0c00082b;
		12'h31f:		data <= 32'h00000000;
		12'h320:		data <= 32'h82100024;
		12'h321:		data <= 32'h2402ffce;
		12'h322:		data <= 32'h12020018;
		12'h323:		data <= 32'h00000000;
		12'h324:		data <= 32'h8e420024;
		12'h325:		data <= 32'h00000000;
		12'h326:		data <= 32'h30420009;
		12'h327:		data <= 32'h10400009;
		12'h328:		data <= 32'h00000000;
		12'h329:		data <= 32'h02001021;
		12'h32a:		data <= 32'h8fbf0020;
		12'h32b:		data <= 32'h8fb3001c;
		12'h32c:		data <= 32'h8fb20018;
		12'h32d:		data <= 32'h8fb10014;
		12'h32e:		data <= 32'h8fb00010;
		12'h32f:		data <= 32'h03e00008;
		12'h330:		data <= 32'h27bd0028;
		12'h331:		data <= 32'h0c00078e;
		12'h332:		data <= 32'h00000000;
		12'h333:		data <= 32'h02001021;
		12'h334:		data <= 32'h8fbf0020;
		12'h335:		data <= 32'h8fb3001c;
		12'h336:		data <= 32'h8fb20018;
		12'h337:		data <= 32'h8fb10014;
		12'h338:		data <= 32'h8fb00010;
		12'h339:		data <= 32'h03e00008;
		12'h33a:		data <= 32'h27bd0028;
		12'h33b:		data <= 32'h08000324;
		12'h33c:		data <= 32'h00008021;
		12'h33d:		data <= 32'h14a0ffeb;
		12'h33e:		data <= 32'h2410ffe7;
		12'h33f:		data <= 32'h0c00078e;
		12'h340:		data <= 32'h00000000;
		12'h341:		data <= 32'h0800032a;
		12'h342:		data <= 32'h02001021;
		12'h343:		data <= 32'h27bdffe0;
		12'h344:		data <= 32'hafb00010;
		12'h345:		data <= 32'hafbf0018;
		12'h346:		data <= 32'hafb10014;
		12'h347:		data <= 32'h1c800007;
		12'h348:		data <= 32'h00808021;
		12'h349:		data <= 32'h2402ffee;
		12'h34a:		data <= 32'h8fbf0018;
		12'h34b:		data <= 32'h8fb10014;
		12'h34c:		data <= 32'h8fb00010;
		12'h34d:		data <= 32'h03e00008;
		12'h34e:		data <= 32'h27bd0020;
		12'h34f:		data <= 32'h3c030000;
		12'h350:		data <= 32'h8c622e90;
		12'h351:		data <= 32'h00000000;
		12'h352:		data <= 32'h0044102a;
		12'h353:		data <= 32'h1440fff6;
		12'h354:		data <= 32'h2402ffee;
		12'h355:		data <= 32'h0c000786;
		12'h356:		data <= 32'h00000000;
		12'h357:		data <= 32'h3c020100;
		12'h358:		data <= 32'h00101880;
		12'h359:		data <= 32'h24420000;
		12'h35a:		data <= 32'h00621821;
		12'h35b:		data <= 32'h8c70fffc;
		12'h35c:		data <= 32'h00000000;
		12'h35d:		data <= 32'h12000030;
		12'h35e:		data <= 32'h3c030100;
		12'h35f:		data <= 32'h0c00090a;
		12'h360:		data <= 32'h02002021;
		12'h361:		data <= 32'h14400014;
		12'h362:		data <= 32'h00408821;
		12'h363:		data <= 32'h8e030004;
		12'h364:		data <= 32'h8e02000c;
		12'h365:		data <= 32'h00000000;
		12'h366:		data <= 32'h0062102b;
		12'h367:		data <= 32'h1040001e;
		12'h368:		data <= 32'h24620001;
		12'h369:		data <= 32'hae020004;
		12'h36a:		data <= 32'h3c030100;
		12'h36b:		data <= 32'h8c6226bc;
		12'h36c:		data <= 32'h00000000;
		12'h36d:		data <= 32'h30420009;
		12'h36e:		data <= 32'h10400003;
		12'h36f:		data <= 32'h00000000;
		12'h370:		data <= 32'h0800034a;
		12'h371:		data <= 32'h00001021;
		12'h372:		data <= 32'h0c00078e;
		12'h373:		data <= 32'h00000000;
		12'h374:		data <= 32'h0800034a;
		12'h375:		data <= 32'h00001021;
		12'h376:		data <= 32'h00021880;
		12'h377:		data <= 32'h3c020100;
		12'h378:		data <= 32'h24420078;
		12'h379:		data <= 32'h00621821;
		12'h37a:		data <= 32'h8c65fffc;
		12'h37b:		data <= 32'h02202021;
		12'h37c:		data <= 32'h0c00087f;
		12'h37d:		data <= 32'ha0a00024;
		12'h37e:		data <= 32'h3c040100;
		12'h37f:		data <= 32'h248426a4;
		12'h380:		data <= 32'h0c0009b9;
		12'h381:		data <= 32'h02202821;
		12'h382:		data <= 32'h0c00082b;
		12'h383:		data <= 32'h00000000;
		12'h384:		data <= 32'h0800036b;
		12'h385:		data <= 32'h3c030100;
		12'h386:		data <= 32'h3c030100;
		12'h387:		data <= 32'h8c6226bc;
		12'h388:		data <= 32'h00000000;
		12'h389:		data <= 32'h30420009;
		12'h38a:		data <= 32'h1040000e;
		12'h38b:		data <= 32'h00000000;
		12'h38c:		data <= 32'h0800034a;
		12'h38d:		data <= 32'h2402ffd5;
		12'h38e:		data <= 32'h8c6226bc;
		12'h38f:		data <= 32'h00000000;
		12'h390:		data <= 32'h30420009;
		12'h391:		data <= 32'h10400003;
		12'h392:		data <= 32'h00000000;
		12'h393:		data <= 32'h0800034a;
		12'h394:		data <= 32'h2402ffd6;
		12'h395:		data <= 32'h0c00078e;
		12'h396:		data <= 32'h00000000;
		12'h397:		data <= 32'h0800034a;
		12'h398:		data <= 32'h2402ffd6;
		12'h399:		data <= 32'h0c00078e;
		12'h39a:		data <= 32'h00000000;
		12'h39b:		data <= 32'h0800034a;
		12'h39c:		data <= 32'h2402ffd5;
		12'h39d:		data <= 32'h080003a1;
		12'h39e:		data <= 32'h2405ffff;
		12'h39f:		data <= 32'h080003a1;
		12'h3a0:		data <= 32'h00002821;
		12'h3a1:		data <= 32'h27bdffd0;
		12'h3a2:		data <= 32'hafb10014;
		12'h3a3:		data <= 32'hafb00010;
		12'h3a4:		data <= 32'hafbf0028;
		12'h3a5:		data <= 32'hafb50024;
		12'h3a6:		data <= 32'hafb40020;
		12'h3a7:		data <= 32'hafb3001c;
		12'h3a8:		data <= 32'hafb20018;
		12'h3a9:		data <= 32'h00a08821;
		12'h3aa:		data <= 32'h10a00006;
		12'h3ab:		data <= 32'h00808021;
		12'h3ac:		data <= 32'h3c020100;
		12'h3ad:		data <= 32'h8c4326bc;
		12'h3ae:		data <= 32'h00000000;
		12'h3af:		data <= 32'h1460000e;
		12'h3b0:		data <= 32'h00000000;
		12'h3b1:		data <= 32'h1e000017;
		12'h3b2:		data <= 32'h3c030000;
		12'h3b3:		data <= 32'h2410ffee;
		12'h3b4:		data <= 32'h02001021;
		12'h3b5:		data <= 32'h8fbf0028;
		12'h3b6:		data <= 32'h8fb50024;
		12'h3b7:		data <= 32'h8fb40020;
		12'h3b8:		data <= 32'h8fb3001c;
		12'h3b9:		data <= 32'h8fb20018;
		12'h3ba:		data <= 32'h8fb10014;
		12'h3bb:		data <= 32'h8fb00010;
		12'h3bc:		data <= 32'h03e00008;
		12'h3bd:		data <= 32'h27bd0030;
		12'h3be:		data <= 32'h2410ffe7;
		12'h3bf:		data <= 32'h02001021;
		12'h3c0:		data <= 32'h8fbf0028;
		12'h3c1:		data <= 32'h8fb50024;
		12'h3c2:		data <= 32'h8fb40020;
		12'h3c3:		data <= 32'h8fb3001c;
		12'h3c4:		data <= 32'h8fb20018;
		12'h3c5:		data <= 32'h8fb10014;
		12'h3c6:		data <= 32'h8fb00010;
		12'h3c7:		data <= 32'h03e00008;
		12'h3c8:		data <= 32'h27bd0030;
		12'h3c9:		data <= 32'h8c622e90;
		12'h3ca:		data <= 32'h00000000;
		12'h3cb:		data <= 32'h0050102a;
		12'h3cc:		data <= 32'h1440ffe6;
		12'h3cd:		data <= 32'h00000000;
		12'h3ce:		data <= 32'h0c000786;
		12'h3cf:		data <= 32'h00000000;
		12'h3d0:		data <= 32'h3c020100;
		12'h3d1:		data <= 32'h00101880;
		12'h3d2:		data <= 32'h24420000;
		12'h3d3:		data <= 32'h00621821;
		12'h3d4:		data <= 32'h8c72fffc;
		12'h3d5:		data <= 32'h00000000;
		12'h3d6:		data <= 32'h12400032;
		12'h3d7:		data <= 32'h3c030100;
		12'h3d8:		data <= 32'h8e420004;
		12'h3d9:		data <= 32'h00000000;
		12'h3da:		data <= 32'h1040000e;
		12'h3db:		data <= 32'h2442ffff;
		12'h3dc:		data <= 32'h00008021;
		12'h3dd:		data <= 32'h3c150100;
		12'h3de:		data <= 32'hae420004;
		12'h3df:		data <= 32'h26a32698;
		12'h3e0:		data <= 32'h8c620024;
		12'h3e1:		data <= 32'h00000000;
		12'h3e2:		data <= 32'h30420009;
		12'h3e3:		data <= 32'h1440ffd0;
		12'h3e4:		data <= 32'h00000000;
		12'h3e5:		data <= 32'h0c00078e;
		12'h3e6:		data <= 32'h00000000;
		12'h3e7:		data <= 32'h080003b5;
		12'h3e8:		data <= 32'h02001021;
		12'h3e9:		data <= 32'h16200003;
		12'h3ea:		data <= 32'h3c150100;
		12'h3eb:		data <= 32'h080003df;
		12'h3ec:		data <= 32'h2410ffce;
		12'h3ed:		data <= 32'h26a22698;
		12'h3ee:		data <= 32'h8c53002c;
		12'h3ef:		data <= 32'h3c020100;
		12'h3f0:		data <= 32'h24420078;
		12'h3f1:		data <= 32'h00131880;
		12'h3f2:		data <= 32'h00621821;
		12'h3f3:		data <= 32'h8c74fffc;
		12'h3f4:		data <= 32'h24020002;
		12'h3f5:		data <= 32'ha282001b;
		12'h3f6:		data <= 32'h02602021;
		12'h3f7:		data <= 32'h0c000874;
		12'h3f8:		data <= 32'ha290001c;
		12'h3f9:		data <= 32'h92460008;
		12'h3fa:		data <= 32'h02402021;
		12'h3fb:		data <= 32'h0c000896;
		12'h3fc:		data <= 32'h02602821;
		12'h3fd:		data <= 32'h2402ffff;
		12'h3fe:		data <= 32'h12220005;
		12'h3ff:		data <= 32'h3c040100;
		12'h400:		data <= 32'h248426a4;
		12'h401:		data <= 32'h02602821;
		12'h402:		data <= 32'h0c000980;
		12'h403:		data <= 32'h02203021;
		12'h404:		data <= 32'h0c00082b;
		12'h405:		data <= 32'h00000000;
		12'h406:		data <= 32'h82900024;
		12'h407:		data <= 32'h080003e0;
		12'h408:		data <= 32'h26a32698;
		12'h409:		data <= 32'h8c6226bc;
		12'h40a:		data <= 32'h00000000;
		12'h40b:		data <= 32'h30420009;
		12'h40c:		data <= 32'h1440ffa7;
		12'h40d:		data <= 32'h2410ffd6;
		12'h40e:		data <= 32'h0c00078e;
		12'h40f:		data <= 32'h00000000;
		12'h410:		data <= 32'h080003b5;
		12'h411:		data <= 32'h02001021;
		12'h412:		data <= 32'h080003a1;
		12'h413:		data <= 32'h00000000;
		12'h414:		data <= 32'h27bdffe0;
		12'h415:		data <= 32'hafb10014;
		12'h416:		data <= 32'hafbf0018;
		12'h417:		data <= 32'h00808821;
		12'h418:		data <= 32'h0c000786;
		12'h419:		data <= 32'hafb00010;
		12'h41a:		data <= 32'h3c020000;
		12'h41b:		data <= 32'h8c442e88;
		12'h41c:		data <= 32'h00000000;
		12'h41d:		data <= 32'h18800032;
		12'h41e:		data <= 32'h3c020100;
		12'h41f:		data <= 32'h2490ffff;
		12'h420:		data <= 32'h24450478;
		12'h421:		data <= 32'h00101880;
		12'h422:		data <= 32'h00651821;
		12'h423:		data <= 32'h8c620000;
		12'h424:		data <= 32'h00000000;
		12'h425:		data <= 32'h10400036;
		12'h426:		data <= 32'h00041080;
		12'h427:		data <= 32'h2442fff8;
		12'h428:		data <= 32'h0800042b;
		12'h429:		data <= 32'h00451821;
		12'h42a:		data <= 32'h00808021;
		12'h42b:		data <= 32'h1a000024;
		12'h42c:		data <= 32'h2604ffff;
		12'h42d:		data <= 32'h8c620000;
		12'h42e:		data <= 32'h00000000;
		12'h42f:		data <= 32'h1440fffa;
		12'h430:		data <= 32'h2463fffc;
		12'h431:		data <= 32'h02202821;
		12'h432:		data <= 32'h0c000462;
		12'h433:		data <= 32'h02002021;
		12'h434:		data <= 32'h1040000d;
		12'h435:		data <= 32'h00408821;
		12'h436:		data <= 32'h3c030100;
		12'h437:		data <= 32'h8c6226bc;
		12'h438:		data <= 32'h00000000;
		12'h439:		data <= 32'h30420009;
		12'h43a:		data <= 32'h1040000d;
		12'h43b:		data <= 32'h00000000;
		12'h43c:		data <= 32'h02201021;
		12'h43d:		data <= 32'h8fbf0018;
		12'h43e:		data <= 32'h8fb10014;
		12'h43f:		data <= 32'h8fb00010;
		12'h440:		data <= 32'h03e00008;
		12'h441:		data <= 32'h27bd0020;
		12'h442:		data <= 32'h3c030100;
		12'h443:		data <= 32'h8c6226bc;
		12'h444:		data <= 32'h00000000;
		12'h445:		data <= 32'h30420009;
		12'h446:		data <= 32'h1440fff5;
		12'h447:		data <= 32'h02008821;
		12'h448:		data <= 32'h0c00078e;
		12'h449:		data <= 32'h00000000;
		12'h44a:		data <= 32'h02201021;
		12'h44b:		data <= 32'h8fbf0018;
		12'h44c:		data <= 32'h8fb10014;
		12'h44d:		data <= 32'h8fb00010;
		12'h44e:		data <= 32'h03e00008;
		12'h44f:		data <= 32'h27bd0020;
		12'h450:		data <= 32'h3c030100;
		12'h451:		data <= 32'h8c6226bc;
		12'h452:		data <= 32'h00000000;
		12'h453:		data <= 32'h30420009;
		12'h454:		data <= 32'h10400009;
		12'h455:		data <= 32'h2411ffde;
		12'h456:		data <= 32'h02201021;
		12'h457:		data <= 32'h8fbf0018;
		12'h458:		data <= 32'h8fb10014;
		12'h459:		data <= 32'h8fb00010;
		12'h45a:		data <= 32'h03e00008;
		12'h45b:		data <= 32'h27bd0020;
		12'h45c:		data <= 32'h08000431;
		12'h45d:		data <= 32'h00808021;
		12'h45e:		data <= 32'h0c00078e;
		12'h45f:		data <= 32'h00000000;
		12'h460:		data <= 32'h08000457;
		12'h461:		data <= 32'h02201021;
		12'h462:		data <= 32'h27bdffe0;
		12'h463:		data <= 32'hafb10014;
		12'h464:		data <= 32'hafb00010;
		12'h465:		data <= 32'hafbf0018;
		12'h466:		data <= 32'h8ca20000;
		12'h467:		data <= 32'h00a08021;
		12'h468:		data <= 32'h30420002;
		12'h469:		data <= 32'h10400005;
		12'h46a:		data <= 32'h00808821;
		12'h46b:		data <= 32'h8ca20008;
		12'h46c:		data <= 32'h00000000;
		12'h46d:		data <= 32'h10400031;
		12'h46e:		data <= 32'h2403ffe0;
		12'h46f:		data <= 32'h24050020;
		12'h470:		data <= 32'h3c040100;
		12'h471:		data <= 32'h0c000a0b;
		12'h472:		data <= 32'h248426b4;
		12'h473:		data <= 32'h10400034;
		12'h474:		data <= 32'h00403021;
		12'h475:		data <= 32'h8e050008;
		12'h476:		data <= 32'h00000000;
		12'h477:		data <= 32'h10a0002e;
		12'h478:		data <= 32'h00000000;
		12'h479:		data <= 32'h3c020100;
		12'h47a:		data <= 32'h8e040000;
		12'h47b:		data <= 32'h24420478;
		12'h47c:		data <= 32'h00111880;
		12'h47d:		data <= 32'h00621821;
		12'h47e:		data <= 32'hac66fffc;
		12'h47f:		data <= 32'ha0c40008;
		12'h480:		data <= 32'h8e030004;
		12'h481:		data <= 32'hacc00000;
		12'h482:		data <= 32'hacc3000c;
		12'h483:		data <= 32'h8e020000;
		12'h484:		data <= 32'h00000000;
		12'h485:		data <= 32'h30420002;
		12'h486:		data <= 32'h10400012;
		12'h487:		data <= 32'h00001021;
		12'h488:		data <= 32'h8e040004;
		12'h489:		data <= 32'h00000000;
		12'h48a:		data <= 32'h18800008;
		12'h48b:		data <= 32'hacc50004;
		12'h48c:		data <= 32'h00a01821;
		12'h48d:		data <= 32'h00003021;
		12'h48e:		data <= 32'h24c60001;
		12'h48f:		data <= 32'h00c4102a;
		12'h490:		data <= 32'hac600000;
		12'h491:		data <= 32'h1440fffc;
		12'h492:		data <= 32'h24630004;
		12'h493:		data <= 32'h8fbf0018;
		12'h494:		data <= 32'h8fb10014;
		12'h495:		data <= 32'h8fb00010;
		12'h496:		data <= 32'h00001021;
		12'h497:		data <= 32'h03e00008;
		12'h498:		data <= 32'h27bd0020;
		12'h499:		data <= 32'hacc00004;
		12'h49a:		data <= 32'h8fbf0018;
		12'h49b:		data <= 32'h8fb10014;
		12'h49c:		data <= 32'h8fb00010;
		12'h49d:		data <= 32'h03e00008;
		12'h49e:		data <= 32'h27bd0020;
		12'h49f:		data <= 32'h8ca20004;
		12'h4a0:		data <= 32'h00000000;
		12'h4a1:		data <= 32'h00021080;
		12'h4a2:		data <= 32'h2442001f;
		12'h4a3:		data <= 32'h00431024;
		12'h4a4:		data <= 32'h08000470;
		12'h4a5:		data <= 32'h24450020;
		12'h4a6:		data <= 32'h08000479;
		12'h4a7:		data <= 32'h24450020;
		12'h4a8:		data <= 32'h8fbf0018;
		12'h4a9:		data <= 32'h8fb10014;
		12'h4aa:		data <= 32'h8fb00010;
		12'h4ab:		data <= 32'h2402ffdf;
		12'h4ac:		data <= 32'h03e00008;
		12'h4ad:		data <= 32'h27bd0020;
		12'h4ae:		data <= 32'h27bdffe0;
		12'h4af:		data <= 32'hafbf001c;
		12'h4b0:		data <= 32'hafb20018;
		12'h4b1:		data <= 32'hafb10014;
		12'h4b2:		data <= 32'hafb00010;
		12'h4b3:		data <= 32'h00a09021;
		12'h4b4:		data <= 32'h0c000786;
		12'h4b5:		data <= 32'h00808021;
		12'h4b6:		data <= 32'h3c020100;
		12'h4b7:		data <= 32'h24420478;
		12'h4b8:		data <= 32'h00108080;
		12'h4b9:		data <= 32'h02028021;
		12'h4ba:		data <= 32'h8e11fffc;
		12'h4bb:		data <= 32'h0c00090a;
		12'h4bc:		data <= 32'h02202021;
		12'h4bd:		data <= 32'h00408021;
		12'h4be:		data <= 32'h00021880;
		12'h4bf:		data <= 32'h3c020100;
		12'h4c0:		data <= 32'h24420078;
		12'h4c1:		data <= 32'h00621821;
		12'h4c2:		data <= 32'h1600001b;
		12'h4c3:		data <= 32'h02002021;
		12'h4c4:		data <= 32'h92220008;
		12'h4c5:		data <= 32'h02202021;
		12'h4c6:		data <= 32'h30420002;
		12'h4c7:		data <= 32'h10400012;
		12'h4c8:		data <= 32'h02402821;
		12'h4c9:		data <= 32'h0c00054e;
		12'h4ca:		data <= 32'h00000000;
		12'h4cb:		data <= 32'h3c030100;
		12'h4cc:		data <= 32'h8c6226bc;
		12'h4cd:		data <= 32'h00000000;
		12'h4ce:		data <= 32'h30420009;
		12'h4cf:		data <= 32'h14400003;
		12'h4d0:		data <= 32'h00000000;
		12'h4d1:		data <= 32'h0c00078e;
		12'h4d2:		data <= 32'h00000000;
		12'h4d3:		data <= 32'h8fbf001c;
		12'h4d4:		data <= 32'h8fb20018;
		12'h4d5:		data <= 32'h8fb10014;
		12'h4d6:		data <= 32'h8fb00010;
		12'h4d7:		data <= 32'h00001021;
		12'h4d8:		data <= 32'h03e00008;
		12'h4d9:		data <= 32'h27bd0020;
		12'h4da:		data <= 32'h0c00054c;
		12'h4db:		data <= 32'h02402821;
		12'h4dc:		data <= 32'h080004cc;
		12'h4dd:		data <= 32'h3c030100;
		12'h4de:		data <= 32'h8c62fffc;
		12'h4df:		data <= 32'h00000000;
		12'h4e0:		data <= 32'h8c430028;
		12'h4e1:		data <= 32'h00000000;
		12'h4e2:		data <= 32'hac720000;
		12'h4e3:		data <= 32'h0c00087f;
		12'h4e4:		data <= 32'ha0400024;
		12'h4e5:		data <= 32'h3c040100;
		12'h4e6:		data <= 32'h248426a4;
		12'h4e7:		data <= 32'h0c0009b9;
		12'h4e8:		data <= 32'h02002821;
		12'h4e9:		data <= 32'h0c00082b;
		12'h4ea:		data <= 32'h00000000;
		12'h4eb:		data <= 32'h080004cc;
		12'h4ec:		data <= 32'h3c030100;
		12'h4ed:		data <= 32'h27bdffd0;
		12'h4ee:		data <= 32'hafb40020;
		12'h4ef:		data <= 32'hafb20018;
		12'h4f0:		data <= 32'hafbf0028;
		12'h4f1:		data <= 32'hafb50024;
		12'h4f2:		data <= 32'hafb3001c;
		12'h4f3:		data <= 32'hafb10014;
		12'h4f4:		data <= 32'hafb00010;
		12'h4f5:		data <= 32'h00809021;
		12'h4f6:		data <= 32'h1c80000c;
		12'h4f7:		data <= 32'h00a0a021;
		12'h4f8:		data <= 32'h2410ffee;
		12'h4f9:		data <= 32'h02001021;
		12'h4fa:		data <= 32'h8fbf0028;
		12'h4fb:		data <= 32'h8fb50024;
		12'h4fc:		data <= 32'h8fb40020;
		12'h4fd:		data <= 32'h8fb3001c;
		12'h4fe:		data <= 32'h8fb20018;
		12'h4ff:		data <= 32'h8fb10014;
		12'h500:		data <= 32'h8fb00010;
		12'h501:		data <= 32'h03e00008;
		12'h502:		data <= 32'h27bd0030;
		12'h503:		data <= 32'h3c030000;
		12'h504:		data <= 32'h8c622e88;
		12'h505:		data <= 32'h00000000;
		12'h506:		data <= 32'h0044102a;
		12'h507:		data <= 32'h1440fff1;
		12'h508:		data <= 32'h2410ffee;
		12'h509:		data <= 32'h0c000786;
		12'h50a:		data <= 32'h00000000;
		12'h50b:		data <= 32'h3c020100;
		12'h50c:		data <= 32'h00121880;
		12'h50d:		data <= 32'h24420478;
		12'h50e:		data <= 32'h00621821;
		12'h50f:		data <= 32'h8c73fffc;
		12'h510:		data <= 32'h00000000;
		12'h511:		data <= 32'h12600031;
		12'h512:		data <= 32'h3c030100;
		12'h513:		data <= 32'h92620008;
		12'h514:		data <= 32'h00000000;
		12'h515:		data <= 32'h30420002;
		12'h516:		data <= 32'h10400012;
		12'h517:		data <= 32'h00000000;
		12'h518:		data <= 32'h8e65000c;
		12'h519:		data <= 32'h0c000569;
		12'h51a:		data <= 32'h02602021;
		12'h51b:		data <= 32'h10400011;
		12'h51c:		data <= 32'h3c150100;
		12'h51d:		data <= 32'h00008021;
		12'h51e:		data <= 32'hae820000;
		12'h51f:		data <= 32'h26a32698;
		12'h520:		data <= 32'h8c620024;
		12'h521:		data <= 32'h00000000;
		12'h522:		data <= 32'h30420009;
		12'h523:		data <= 32'h1440ffd5;
		12'h524:		data <= 32'h00000000;
		12'h525:		data <= 32'h0c00078e;
		12'h526:		data <= 32'h00000000;
		12'h527:		data <= 32'h080004fa;
		12'h528:		data <= 32'h02001021;
		12'h529:		data <= 32'h0c000561;
		12'h52a:		data <= 32'h02602021;
		12'h52b:		data <= 32'h0800051b;
		12'h52c:		data <= 32'h00000000;
		12'h52d:		data <= 32'h26a22698;
		12'h52e:		data <= 32'h8c51002c;
		12'h52f:		data <= 32'h3c020100;
		12'h530:		data <= 32'h24420078;
		12'h531:		data <= 32'h00111880;
		12'h532:		data <= 32'h00621821;
		12'h533:		data <= 32'h8c70fffc;
		12'h534:		data <= 32'h24020002;
		12'h535:		data <= 32'ha202001b;
		12'h536:		data <= 32'ha212001c;
		12'h537:		data <= 32'hae140028;
		12'h538:		data <= 32'h0c000874;
		12'h539:		data <= 32'h02202021;
		12'h53a:		data <= 32'h92660008;
		12'h53b:		data <= 32'h02602021;
		12'h53c:		data <= 32'h0c000896;
		12'h53d:		data <= 32'h02202821;
		12'h53e:		data <= 32'h0c00082b;
		12'h53f:		data <= 32'h00000000;
		12'h540:		data <= 32'h82100024;
		12'h541:		data <= 32'h08000520;
		12'h542:		data <= 32'h26a32698;
		12'h543:		data <= 32'h8c6226bc;
		12'h544:		data <= 32'h00000000;
		12'h545:		data <= 32'h30420009;
		12'h546:		data <= 32'h1440ffb2;
		12'h547:		data <= 32'h2410ffd6;
		12'h548:		data <= 32'h0c00078e;
		12'h549:		data <= 32'h00000000;
		12'h54a:		data <= 32'h080004fa;
		12'h54b:		data <= 32'h02001021;
		12'h54c:		data <= 32'h08000554;
		12'h54d:		data <= 32'h24840004;
		12'h54e:		data <= 32'h8ca20004;
		12'h54f:		data <= 32'h8c840004;
		12'h550:		data <= 32'h00021080;
		12'h551:		data <= 32'h00822021;
		12'h552:		data <= 32'h08000554;
		12'h553:		data <= 32'h2484fffc;
		12'h554:		data <= 32'h8c830000;
		12'h555:		data <= 32'h00000000;
		12'h556:		data <= 32'h10600007;
		12'h557:		data <= 32'h00000000;
		12'h558:		data <= 32'h8c620000;
		12'h559:		data <= 32'h00000000;
		12'h55a:		data <= 32'haca20000;
		12'h55b:		data <= 32'hac650000;
		12'h55c:		data <= 32'h03e00008;
		12'h55d:		data <= 32'hac850000;
		12'h55e:		data <= 32'haca50000;
		12'h55f:		data <= 32'h03e00008;
		12'h560:		data <= 32'hac850000;
		12'h561:		data <= 32'h8c820004;
		12'h562:		data <= 32'h00000000;
		12'h563:		data <= 32'h10400003;
		12'h564:		data <= 32'h24840004;
		12'h565:		data <= 32'h08000582;
		12'h566:		data <= 32'h00000000;
		12'h567:		data <= 32'h03e00008;
		12'h568:		data <= 32'h00001021;
		12'h569:		data <= 32'h28a20002;
		12'h56a:		data <= 32'h14400009;
		12'h56b:		data <= 32'h00000000;
		12'h56c:		data <= 32'h8c840004;
		12'h56d:		data <= 32'h00000000;
		12'h56e:		data <= 32'h8c820004;
		12'h56f:		data <= 32'h00000000;
		12'h570:		data <= 32'h10400005;
		12'h571:		data <= 32'h24830004;
		12'h572:		data <= 32'h08000582;
		12'h573:		data <= 32'h00602021;
		12'h574:		data <= 32'h03e00008;
		12'h575:		data <= 32'h00001021;
		12'h576:		data <= 32'h24840008;
		12'h577:		data <= 32'h24060001;
		12'h578:		data <= 32'h24c60001;
		12'h579:		data <= 32'h00801821;
		12'h57a:		data <= 32'h10a6fff9;
		12'h57b:		data <= 32'h24840004;
		12'h57c:		data <= 32'h8c620000;
		12'h57d:		data <= 32'h00000000;
		12'h57e:		data <= 32'h1040fffa;
		12'h57f:		data <= 32'h24c60001;
		12'h580:		data <= 32'h08000582;
		12'h581:		data <= 32'h00602021;
		12'h582:		data <= 32'h8c830000;
		12'h583:		data <= 32'h00000000;
		12'h584:		data <= 32'h8c650000;
		12'h585:		data <= 32'h00000000;
		12'h586:		data <= 32'h10650006;
		12'h587:		data <= 32'h00000000;
		12'h588:		data <= 32'h8ca20000;
		12'h589:		data <= 32'h00000000;
		12'h58a:		data <= 32'hac620000;
		12'h58b:		data <= 32'h03e00008;
		12'h58c:		data <= 32'h00a01021;
		12'h58d:		data <= 32'h00a01021;
		12'h58e:		data <= 32'h03e00008;
		12'h58f:		data <= 32'hac800000;
		12'h590:		data <= 32'h27bdffe0;
		12'h591:		data <= 32'hafb10014;
		12'h592:		data <= 32'hafbf0018;
		12'h593:		data <= 32'hafb00010;
		12'h594:		data <= 32'h0c000786;
		12'h595:		data <= 32'h00808821;
		12'h596:		data <= 32'h3c020000;
		12'h597:		data <= 32'h8c452e80;
		12'h598:		data <= 32'h00000000;
		12'h599:		data <= 32'h18a0002a;
		12'h59a:		data <= 32'h24b0ffff;
		12'h59b:		data <= 32'h001020c0;
		12'h59c:		data <= 32'h3c030100;
		12'h59d:		data <= 32'h00101140;
		12'h59e:		data <= 32'h00441023;
		12'h59f:		data <= 32'h2464024c;
		12'h5a0:		data <= 32'h00441021;
		12'h5a1:		data <= 32'h8c430014;
		12'h5a2:		data <= 32'h00000000;
		12'h5a3:		data <= 32'h1060002c;
		12'h5a4:		data <= 32'h000518c0;
		12'h5a5:		data <= 32'h00051140;
		12'h5a6:		data <= 32'h00431023;
		12'h5a7:		data <= 32'h00441021;
		12'h5a8:		data <= 32'h080005ab;
		12'h5a9:		data <= 32'h2443ffe4;
		12'h5aa:		data <= 32'h00808021;
		12'h5ab:		data <= 32'h1a000018;
		12'h5ac:		data <= 32'h2604ffff;
		12'h5ad:		data <= 32'h8c620000;
		12'h5ae:		data <= 32'h00000000;
		12'h5af:		data <= 32'h1440fffa;
		12'h5b0:		data <= 32'h2463ffe8;
		12'h5b1:		data <= 32'h02202821;
		12'h5b2:		data <= 32'h0c0005e1;
		12'h5b3:		data <= 32'h02002021;
		12'h5b4:		data <= 32'h3c030100;
		12'h5b5:		data <= 32'h8c6226bc;
		12'h5b6:		data <= 32'h00000000;
		12'h5b7:		data <= 32'h30420009;
		12'h5b8:		data <= 32'h10400007;
		12'h5b9:		data <= 32'h00000000;
		12'h5ba:		data <= 32'h02001021;
		12'h5bb:		data <= 32'h8fbf0018;
		12'h5bc:		data <= 32'h8fb10014;
		12'h5bd:		data <= 32'h8fb00010;
		12'h5be:		data <= 32'h03e00008;
		12'h5bf:		data <= 32'h27bd0020;
		12'h5c0:		data <= 32'h0c00078e;
		12'h5c1:		data <= 32'h00000000;
		12'h5c2:		data <= 32'h080005bb;
		12'h5c3:		data <= 32'h02001021;
		12'h5c4:		data <= 32'h3c030100;
		12'h5c5:		data <= 32'h8c6226bc;
		12'h5c6:		data <= 32'h00000000;
		12'h5c7:		data <= 32'h30420009;
		12'h5c8:		data <= 32'h10400009;
		12'h5c9:		data <= 32'h00000000;
		12'h5ca:		data <= 32'h2402ffde;
		12'h5cb:		data <= 32'h8fbf0018;
		12'h5cc:		data <= 32'h8fb10014;
		12'h5cd:		data <= 32'h8fb00010;
		12'h5ce:		data <= 32'h03e00008;
		12'h5cf:		data <= 32'h27bd0020;
		12'h5d0:		data <= 32'h080005b1;
		12'h5d1:		data <= 32'h00a08021;
		12'h5d2:		data <= 32'h0c00078e;
		12'h5d3:		data <= 32'h00000000;
		12'h5d4:		data <= 32'h080005cb;
		12'h5d5:		data <= 32'h2402ffde;
		12'h5d6:		data <= 32'h24a5ffff;
		12'h5d7:		data <= 32'h24020001;
		12'h5d8:		data <= 32'h2ca30002;
		12'h5d9:		data <= 32'h14600005;
		12'h5da:		data <= 32'hac820004;
		12'h5db:		data <= 32'h24420001;
		12'h5dc:		data <= 32'hace20000;
		12'h5dd:		data <= 32'h1445fffd;
		12'h5de:		data <= 32'h00e63821;
		12'h5df:		data <= 32'h03e00008;
		12'h5e0:		data <= 32'hace00000;
		12'h5e1:		data <= 32'h27bdffe0;
		12'h5e2:		data <= 32'hafb10014;
		12'h5e3:		data <= 32'hafb00010;
		12'h5e4:		data <= 32'hafbf0018;
		12'h5e5:		data <= 32'h8caa000c;
		12'h5e6:		data <= 32'h00808821;
		12'h5e7:		data <= 32'h3c040100;
		12'h5e8:		data <= 32'h00a08021;
		12'h5e9:		data <= 32'h1140001e;
		12'h5ea:		data <= 32'h248426b4;
		12'h5eb:		data <= 32'h001110c0;
		12'h5ec:		data <= 32'h00111940;
		12'h5ed:		data <= 32'h00621823;
		12'h5ee:		data <= 32'h3c020100;
		12'h5ef:		data <= 32'h2442024c;
		12'h5f0:		data <= 32'h8e040000;
		12'h5f1:		data <= 32'h2442ffe8;
		12'h5f2:		data <= 32'h00621821;
		12'h5f3:		data <= 32'ha0640008;
		12'h5f4:		data <= 32'h8e080008;
		12'h5f5:		data <= 32'h8e090004;
		12'h5f6:		data <= 32'h2402fffc;
		12'h5f7:		data <= 32'hac600000;
		12'h5f8:		data <= 32'h25080003;
		12'h5f9:		data <= 32'h01024024;
		12'h5fa:		data <= 32'h8e060008;
		12'h5fb:		data <= 32'h8e050004;
		12'h5fc:		data <= 32'h00602021;
		12'h5fd:		data <= 32'h01403821;
		12'h5fe:		data <= 32'hac69000c;
		12'h5ff:		data <= 32'hac680010;
		12'h600:		data <= 32'h0c0005d6;
		12'h601:		data <= 32'hac6a0014;
		12'h602:		data <= 32'h00001021;
		12'h603:		data <= 32'h8fbf0018;
		12'h604:		data <= 32'h8fb10014;
		12'h605:		data <= 32'h8fb00010;
		12'h606:		data <= 32'h03e00008;
		12'h607:		data <= 32'h27bd0020;
		12'h608:		data <= 32'h8ca50008;
		12'h609:		data <= 32'h8e030004;
		12'h60a:		data <= 32'h2402fffc;
		12'h60b:		data <= 32'h24a50003;
		12'h60c:		data <= 32'h00a22824;
		12'h60d:		data <= 32'h00650018;
		12'h60e:		data <= 32'h00002812;
		12'h60f:		data <= 32'h0c000a0b;
		12'h610:		data <= 32'h00000000;
		12'h611:		data <= 32'h00405021;
		12'h612:		data <= 32'h1540ffd8;
		12'h613:		data <= 32'h2402ffdf;
		12'h614:		data <= 32'h08000603;
		12'h615:		data <= 32'h00000000;
		12'h616:		data <= 32'h27bdffd0;
		12'h617:		data <= 32'hafb3001c;
		12'h618:		data <= 32'h3c130100;
		12'h619:		data <= 32'hafb40020;
		12'h61a:		data <= 32'hafb20018;
		12'h61b:		data <= 32'hafb00010;
		12'h61c:		data <= 32'hafbf0028;
		12'h61d:		data <= 32'hafb50024;
		12'h61e:		data <= 32'hafb10014;
		12'h61f:		data <= 32'h26702698;
		12'h620:		data <= 32'h8e020024;
		12'h621:		data <= 32'h00809021;
		12'h622:		data <= 32'h1040000c;
		12'h623:		data <= 32'h00a0a021;
		12'h624:		data <= 32'h2410ffe7;
		12'h625:		data <= 32'h02001021;
		12'h626:		data <= 32'h8fbf0028;
		12'h627:		data <= 32'h8fb50024;
		12'h628:		data <= 32'h8fb40020;
		12'h629:		data <= 32'h8fb3001c;
		12'h62a:		data <= 32'h8fb20018;
		12'h62b:		data <= 32'h8fb10014;
		12'h62c:		data <= 32'h8fb00010;
		12'h62d:		data <= 32'h03e00008;
		12'h62e:		data <= 32'h27bd0030;
		12'h62f:		data <= 32'h1c800003;
		12'h630:		data <= 32'h3c030000;
		12'h631:		data <= 32'h08000625;
		12'h632:		data <= 32'h2410ffee;
		12'h633:		data <= 32'h8c622e80;
		12'h634:		data <= 32'h00000000;
		12'h635:		data <= 32'h0044102a;
		12'h636:		data <= 32'h1440fffa;
		12'h637:		data <= 32'h00000000;
		12'h638:		data <= 32'h0c000786;
		12'h639:		data <= 32'h00000000;
		12'h63a:		data <= 32'h00121140;
		12'h63b:		data <= 32'h3c030100;
		12'h63c:		data <= 32'h001220c0;
		12'h63d:		data <= 32'h2465024c;
		12'h63e:		data <= 32'h00442023;
		12'h63f:		data <= 32'h00851021;
		12'h640:		data <= 32'h8c43fffc;
		12'h641:		data <= 32'h00000000;
		12'h642:		data <= 32'h1060002e;
		12'h643:		data <= 32'h24a2ffe8;
		12'h644:		data <= 32'h0082a821;
		12'h645:		data <= 32'h8ea30004;
		12'h646:		data <= 32'h00000000;
		12'h647:		data <= 32'h10600015;
		12'h648:		data <= 32'h3c020100;
		12'h649:		data <= 32'h8ea40010;
		12'h64a:		data <= 32'h2463ffff;
		12'h64b:		data <= 32'h00640018;
		12'h64c:		data <= 32'h8ea20014;
		12'h64d:		data <= 32'h00008021;
		12'h64e:		data <= 32'h00001812;
		12'h64f:		data <= 32'h00431021;
		12'h650:		data <= 32'h8c440000;
		12'h651:		data <= 32'hae820000;
		12'h652:		data <= 32'haea40004;
		12'h653:		data <= 32'h26632698;
		12'h654:		data <= 32'h8c620024;
		12'h655:		data <= 32'h00000000;
		12'h656:		data <= 32'h30420009;
		12'h657:		data <= 32'h1440ffcd;
		12'h658:		data <= 32'h00000000;
		12'h659:		data <= 32'h0c00078e;
		12'h65a:		data <= 32'h00000000;
		12'h65b:		data <= 32'h08000626;
		12'h65c:		data <= 32'h02001021;
		12'h65d:		data <= 32'h8e11002c;
		12'h65e:		data <= 32'h24420078;
		12'h65f:		data <= 32'h00111880;
		12'h660:		data <= 32'h00621821;
		12'h661:		data <= 32'h8c70fffc;
		12'h662:		data <= 32'h2402000d;
		12'h663:		data <= 32'ha202001b;
		12'h664:		data <= 32'ha212001c;
		12'h665:		data <= 32'hae140028;
		12'h666:		data <= 32'h0c000874;
		12'h667:		data <= 32'h02202021;
		12'h668:		data <= 32'h92a60008;
		12'h669:		data <= 32'h02a02021;
		12'h66a:		data <= 32'h0c000896;
		12'h66b:		data <= 32'h02202821;
		12'h66c:		data <= 32'h0c00082b;
		12'h66d:		data <= 32'h00000000;
		12'h66e:		data <= 32'h82100024;
		12'h66f:		data <= 32'h08000654;
		12'h670:		data <= 32'h26632698;
		12'h671:		data <= 32'h8e020024;
		12'h672:		data <= 32'h00000000;
		12'h673:		data <= 32'h30420009;
		12'h674:		data <= 32'h14400003;
		12'h675:		data <= 32'h00000000;
		12'h676:		data <= 32'h0c00078e;
		12'h677:		data <= 32'h00000000;
		12'h678:		data <= 32'h08000625;
		12'h679:		data <= 32'h2410ffd6;
		12'h67a:		data <= 32'h27bdffd8;
		12'h67b:		data <= 32'hafb3001c;
		12'h67c:		data <= 32'h3c130100;
		12'h67d:		data <= 32'hafb20018;
		12'h67e:		data <= 32'hafb10014;
		12'h67f:		data <= 32'hafb00010;
		12'h680:		data <= 32'hafbf0020;
		12'h681:		data <= 32'h26712698;
		12'h682:		data <= 32'h8e220024;
		12'h683:		data <= 32'h00808021;
		12'h684:		data <= 32'h1040000c;
		12'h685:		data <= 32'h00a09021;
		12'h686:		data <= 32'h30420009;
		12'h687:		data <= 32'h10400041;
		12'h688:		data <= 32'h00000000;
		12'h689:		data <= 32'h2402ffe7;
		12'h68a:		data <= 32'h8fbf0020;
		12'h68b:		data <= 32'h8fb3001c;
		12'h68c:		data <= 32'h8fb20018;
		12'h68d:		data <= 32'h8fb10014;
		12'h68e:		data <= 32'h8fb00010;
		12'h68f:		data <= 32'h03e00008;
		12'h690:		data <= 32'h27bd0028;
		12'h691:		data <= 32'h1c800009;
		12'h692:		data <= 32'h3c030000;
		12'h693:		data <= 32'h8fbf0020;
		12'h694:		data <= 32'h8fb3001c;
		12'h695:		data <= 32'h8fb20018;
		12'h696:		data <= 32'h8fb10014;
		12'h697:		data <= 32'h8fb00010;
		12'h698:		data <= 32'h2402ffee;
		12'h699:		data <= 32'h03e00008;
		12'h69a:		data <= 32'h27bd0028;
		12'h69b:		data <= 32'h8c622e80;
		12'h69c:		data <= 32'h00000000;
		12'h69d:		data <= 32'h0044102a;
		12'h69e:		data <= 32'h1440fff4;
		12'h69f:		data <= 32'h00000000;
		12'h6a0:		data <= 32'h0c000786;
		12'h6a1:		data <= 32'h00000000;
		12'h6a2:		data <= 32'h001010c0;
		12'h6a3:		data <= 32'h3c030100;
		12'h6a4:		data <= 32'h00102140;
		12'h6a5:		data <= 32'h2465024c;
		12'h6a6:		data <= 32'h00822023;
		12'h6a7:		data <= 32'h00851021;
		12'h6a8:		data <= 32'h8c43fffc;
		12'h6a9:		data <= 32'h00000000;
		12'h6aa:		data <= 32'h10600031;
		12'h6ab:		data <= 32'h24a2ffe8;
		12'h6ac:		data <= 32'h00828021;
		12'h6ad:		data <= 32'h0c00090a;
		12'h6ae:		data <= 32'h02002021;
		12'h6af:		data <= 32'h1440001d;
		12'h6b0:		data <= 32'h00402021;
		12'h6b1:		data <= 32'h8e020014;
		12'h6b2:		data <= 32'h8e040010;
		12'h6b3:		data <= 32'h02421023;
		12'h6b4:		data <= 32'h14800002;
		12'h6b5:		data <= 32'h0044001b;
		12'h6b6:		data <= 32'h0007000d;
		12'h6b7:		data <= 32'h8e030004;
		12'h6b8:		data <= 32'h00000000;
		12'h6b9:		data <= 32'hae430000;
		12'h6ba:		data <= 32'h00001012;
		12'h6bb:		data <= 32'h24420001;
		12'h6bc:		data <= 32'hae020004;
		12'h6bd:		data <= 32'h26632698;
		12'h6be:		data <= 32'h8c620024;
		12'h6bf:		data <= 32'h00000000;
		12'h6c0:		data <= 32'h30420009;
		12'h6c1:		data <= 32'h10400003;
		12'h6c2:		data <= 32'h00000000;
		12'h6c3:		data <= 32'h0800068a;
		12'h6c4:		data <= 32'h00001021;
		12'h6c5:		data <= 32'h0c00078e;
		12'h6c6:		data <= 32'h00000000;
		12'h6c7:		data <= 32'h0800068a;
		12'h6c8:		data <= 32'h00001021;
		12'h6c9:		data <= 32'h0c00078e;
		12'h6ca:		data <= 32'h00000000;
		12'h6cb:		data <= 32'h0800068a;
		12'h6cc:		data <= 32'h2402ffe7;
		12'h6cd:		data <= 32'h00021880;
		12'h6ce:		data <= 32'h3c020100;
		12'h6cf:		data <= 32'h24420078;
		12'h6d0:		data <= 32'h00621821;
		12'h6d1:		data <= 32'h8c65fffc;
		12'h6d2:		data <= 32'h00000000;
		12'h6d3:		data <= 32'h8ca20028;
		12'h6d4:		data <= 32'h00000000;
		12'h6d5:		data <= 32'hac520000;
		12'h6d6:		data <= 32'h0c00087f;
		12'h6d7:		data <= 32'ha0a00024;
		12'h6d8:		data <= 32'h0c00082b;
		12'h6d9:		data <= 32'h00000000;
		12'h6da:		data <= 32'h080006be;
		12'h6db:		data <= 32'h26632698;
		12'h6dc:		data <= 32'h8e220024;
		12'h6dd:		data <= 32'h00000000;
		12'h6de:		data <= 32'h30420009;
		12'h6df:		data <= 32'h10400003;
		12'h6e0:		data <= 32'h00000000;
		12'h6e1:		data <= 32'h0800068a;
		12'h6e2:		data <= 32'h2402ffd6;
		12'h6e3:		data <= 32'h0c00078e;
		12'h6e4:		data <= 32'h00000000;
		12'h6e5:		data <= 32'h0800068a;
		12'h6e6:		data <= 32'h2402ffd6;
		12'h6e7:		data <= 32'h27bdffe8;
		12'h6e8:		data <= 32'hafbf0014;
		12'h6e9:		data <= 32'h0c000786;
		12'h6ea:		data <= 32'hafb00010;
		12'h6eb:		data <= 32'h3c040100;
		12'h6ec:		data <= 32'h3c050000;
		12'h6ed:		data <= 32'h2484269c;
		12'h6ee:		data <= 32'h0c000922;
		12'h6ef:		data <= 32'h24a52e74;
		12'h6f0:		data <= 32'h3c040100;
		12'h6f1:		data <= 32'h00402821;
		12'h6f2:		data <= 32'h248426a8;
		12'h6f3:		data <= 32'h0c0009e0;
		12'h6f4:		data <= 32'h00408021;
		12'h6f5:		data <= 32'h3c040100;
		12'h6f6:		data <= 32'h248426a4;
		12'h6f7:		data <= 32'h0c000940;
		12'h6f8:		data <= 32'h02002821;
		12'h6f9:		data <= 32'h3c030100;
		12'h6fa:		data <= 32'h8c6226bc;
		12'h6fb:		data <= 32'h00000000;
		12'h6fc:		data <= 32'h30420009;
		12'h6fd:		data <= 32'h14400003;
		12'h6fe:		data <= 32'h00000000;
		12'h6ff:		data <= 32'h0c00078e;
		12'h700:		data <= 32'h00000000;
		12'h701:		data <= 32'h8fbf0014;
		12'h702:		data <= 32'h8fb00010;
		12'h703:		data <= 32'h00001021;
		12'h704:		data <= 32'h03e00008;
		12'h705:		data <= 32'h27bd0018;
		12'h706:		data <= 32'h27bdffe0;
		12'h707:		data <= 32'hafb10014;
		12'h708:		data <= 32'hafb00010;
		12'h709:		data <= 32'hafbf0018;
		12'h70a:		data <= 32'h0c000786;
		12'h70b:		data <= 32'h00808821;
		12'h70c:		data <= 32'h3c020000;
		12'h70d:		data <= 32'h8c502e64;
		12'h70e:		data <= 32'h00000000;
		12'h70f:		data <= 32'h1a000014;
		12'h710:		data <= 32'h3c020100;
		12'h711:		data <= 32'h2605ffff;
		12'h712:		data <= 32'h24441688;
		12'h713:		data <= 32'h00051880;
		12'h714:		data <= 32'h00641821;
		12'h715:		data <= 32'h8c620000;
		12'h716:		data <= 32'h00000000;
		12'h717:		data <= 32'h1040000c;
		12'h718:		data <= 32'h00101080;
		12'h719:		data <= 32'h2442fff8;
		12'h71a:		data <= 32'h00442021;
		12'h71b:		data <= 32'h0800071e;
		12'h71c:		data <= 32'h00a08021;
		12'h71d:		data <= 32'h00608021;
		12'h71e:		data <= 32'h1a000026;
		12'h71f:		data <= 32'h2603ffff;
		12'h720:		data <= 32'h8c820000;
		12'h721:		data <= 32'h00000000;
		12'h722:		data <= 32'h1440fffa;
		12'h723:		data <= 32'h2484fffc;
		12'h724:		data <= 32'h2a020002;
		12'h725:		data <= 32'h1440001f;
		12'h726:		data <= 32'h02202821;
		12'h727:		data <= 32'h0c000755;
		12'h728:		data <= 32'h02002021;
		12'h729:		data <= 32'h1040000d;
		12'h72a:		data <= 32'h00408821;
		12'h72b:		data <= 32'h3c030100;
		12'h72c:		data <= 32'h8c6226bc;
		12'h72d:		data <= 32'h00000000;
		12'h72e:		data <= 32'h30420009;
		12'h72f:		data <= 32'h1040000d;
		12'h730:		data <= 32'h00000000;
		12'h731:		data <= 32'h02201021;
		12'h732:		data <= 32'h8fbf0018;
		12'h733:		data <= 32'h8fb10014;
		12'h734:		data <= 32'h8fb00010;
		12'h735:		data <= 32'h03e00008;
		12'h736:		data <= 32'h27bd0020;
		12'h737:		data <= 32'h3c030100;
		12'h738:		data <= 32'h8c6226bc;
		12'h739:		data <= 32'h00000000;
		12'h73a:		data <= 32'h30420009;
		12'h73b:		data <= 32'h1440fff5;
		12'h73c:		data <= 32'h02008821;
		12'h73d:		data <= 32'h0c00078e;
		12'h73e:		data <= 32'h00000000;
		12'h73f:		data <= 32'h02201021;
		12'h740:		data <= 32'h8fbf0018;
		12'h741:		data <= 32'h8fb10014;
		12'h742:		data <= 32'h8fb00010;
		12'h743:		data <= 32'h03e00008;
		12'h744:		data <= 32'h27bd0020;
		12'h745:		data <= 32'h3c030100;
		12'h746:		data <= 32'h8c6226bc;
		12'h747:		data <= 32'h00000000;
		12'h748:		data <= 32'h30420009;
		12'h749:		data <= 32'h10400007;
		12'h74a:		data <= 32'h2411ffde;
		12'h74b:		data <= 32'h02201021;
		12'h74c:		data <= 32'h8fbf0018;
		12'h74d:		data <= 32'h8fb10014;
		12'h74e:		data <= 32'h8fb00010;
		12'h74f:		data <= 32'h03e00008;
		12'h750:		data <= 32'h27bd0020;
		12'h751:		data <= 32'h0c00078e;
		12'h752:		data <= 32'h00000000;
		12'h753:		data <= 32'h0800074c;
		12'h754:		data <= 32'h02201021;
		12'h755:		data <= 32'h27bdffe0;
		12'h756:		data <= 32'hafb20018;
		12'h757:		data <= 32'hafb10014;
		12'h758:		data <= 32'hafb00010;
		12'h759:		data <= 32'h3c020000;
		12'h75a:		data <= 32'hafbf001c;
		12'h75b:		data <= 32'h8c512e6c;
		12'h75c:		data <= 32'h8ca60008;
		12'h75d:		data <= 32'h00a08021;
		12'h75e:		data <= 32'h00d1102a;
		12'h75f:		data <= 32'h10400009;
		12'h760:		data <= 32'h00809021;
		12'h761:		data <= 32'h2403ffef;
		12'h762:		data <= 32'h8fbf001c;
		12'h763:		data <= 32'h8fb20018;
		12'h764:		data <= 32'h8fb10014;
		12'h765:		data <= 32'h8fb00010;
		12'h766:		data <= 32'h00601021;
		12'h767:		data <= 32'h03e00008;
		12'h768:		data <= 32'h27bd0020;
		12'h769:		data <= 32'h3c020000;
		12'h76a:		data <= 32'h8c432e68;
		12'h76b:		data <= 32'h3c040100;
		12'h76c:		data <= 32'h0066182a;
		12'h76d:		data <= 32'h248426b4;
		12'h76e:		data <= 32'h1460fff2;
		12'h76f:		data <= 32'h2405000c;
		12'h770:		data <= 32'h0c000a0b;
		12'h771:		data <= 32'h00000000;
		12'h772:		data <= 32'h8e030004;
		12'h773:		data <= 32'h00122880;
		12'h774:		data <= 32'hac430004;
		12'h775:		data <= 32'h8e040008;
		12'h776:		data <= 32'h3c030100;
		12'h777:		data <= 32'h00912023;
		12'h778:		data <= 32'h24631288;
		12'h779:		data <= 32'h00042080;
		12'h77a:		data <= 32'h00832021;
		12'h77b:		data <= 32'h3c030100;
		12'h77c:		data <= 32'h8c870000;
		12'h77d:		data <= 32'h24631688;
		12'h77e:		data <= 32'h8e06000c;
		12'h77f:		data <= 32'h00a32821;
		12'h780:		data <= 32'h00001821;
		12'h781:		data <= 32'haca2fffc;
		12'h782:		data <= 32'hac460008;
		12'h783:		data <= 32'hac470000;
		12'h784:		data <= 32'h08000762;
		12'h785:		data <= 32'hac820000;
		12'h786:		data <= 32'h40086000;
		12'h787:		data <= 32'h3c09f1ff;
		12'h788:		data <= 32'h3529fff8;
		12'h789:		data <= 32'h01094024;
		12'h78a:		data <= 32'h40886000;
		12'h78b:		data <= 32'h00000000;
		12'h78c:		data <= 32'h03e00008;
		12'h78d:		data <= 32'h00000000;
		12'h78e:		data <= 32'h40086000;
		12'h78f:		data <= 32'h3c09f1ff;
		12'h790:		data <= 32'h3529fffb;
		12'h791:		data <= 32'h01094024;
		12'h792:		data <= 32'h35080001;
		12'h793:		data <= 32'h40886000;
		12'h794:		data <= 32'h00000000;
		12'h795:		data <= 32'h03e00008;
		12'h796:		data <= 32'h00000000;
		12'h797:		data <= 32'h24a5ffd8;
		12'h798:		data <= 32'hac850000;
		12'h799:		data <= 32'h8fa80010;
		12'h79a:		data <= 32'haca70000;
		12'h79b:		data <= 32'haca80004;
		12'h79c:		data <= 32'haca60008;
		12'h79d:		data <= 32'h3c080000;
		12'h79e:		data <= 32'h25081e84;
		12'h79f:		data <= 32'h03e00008;
		12'h7a0:		data <= 32'haca80024;
		12'h7a1:		data <= 32'h02002021;
		12'h7a2:		data <= 32'h02400008;
		12'h7a3:		data <= 32'h02202821;
		12'h7a4:		data <= 32'h27bdffd8;
		12'h7a5:		data <= 32'hafb00000;
		12'h7a6:		data <= 32'hafb10004;
		12'h7a7:		data <= 32'hafb20008;
		12'h7a8:		data <= 32'hafb3000c;
		12'h7a9:		data <= 32'hafb40010;
		12'h7aa:		data <= 32'hafb50014;
		12'h7ab:		data <= 32'hafb60018;
		12'h7ac:		data <= 32'hafb7001c;
		12'h7ad:		data <= 32'hafbe0020;
		12'h7ae:		data <= 32'hafbf0024;
		12'h7af:		data <= 32'hacbd0000;
		12'h7b0:		data <= 32'h8c9d0000;
		12'h7b1:		data <= 32'h00000000;
		12'h7b2:		data <= 32'h8fbf0024;
		12'h7b3:		data <= 32'h8fbe0020;
		12'h7b4:		data <= 32'h8fb7001c;
		12'h7b5:		data <= 32'h8fb60018;
		12'h7b6:		data <= 32'h8fb50014;
		12'h7b7:		data <= 32'h8fb40010;
		12'h7b8:		data <= 32'h8fb3000c;
		12'h7b9:		data <= 32'h8fb20008;
		12'h7ba:		data <= 32'h8fb10004;
		12'h7bb:		data <= 32'h8fb00000;
		12'h7bc:		data <= 32'h03e00008;
		12'h7bd:		data <= 32'h27bd0028;
		12'h7be:		data <= 32'h27bdffac;
		12'h7bf:		data <= 32'hafa10000;
		12'h7c0:		data <= 32'hafa20004;
		12'h7c1:		data <= 32'hafa30008;
		12'h7c2:		data <= 32'hafa4000c;
		12'h7c3:		data <= 32'hafa50010;
		12'h7c4:		data <= 32'hafa60014;
		12'h7c5:		data <= 32'hafa70018;
		12'h7c6:		data <= 32'hafa8001c;
		12'h7c7:		data <= 32'hafa90020;
		12'h7c8:		data <= 32'hafaa0024;
		12'h7c9:		data <= 32'hafab0028;
		12'h7ca:		data <= 32'hafac002c;
		12'h7cb:		data <= 32'hafad0030;
		12'h7cc:		data <= 32'hafae0034;
		12'h7cd:		data <= 32'hafaf0038;
		12'h7ce:		data <= 32'hafb8003c;
		12'h7cf:		data <= 32'hafb90040;
		12'h7d0:		data <= 32'hafbf0044;
		12'h7d1:		data <= 32'h00004010;
		12'h7d2:		data <= 32'h00004812;
		12'h7d3:		data <= 32'h400a7000;
		12'h7d4:		data <= 32'hafa80048;
		12'h7d5:		data <= 32'hafa9004c;
		12'h7d6:		data <= 32'hafaa0050;
		12'h7d7:		data <= 32'h0c000b01;
		12'h7d8:		data <= 32'hafaa004c;
		12'h7d9:		data <= 32'h24040000;
		12'h7da:		data <= 32'h0c000b08;
		12'h7db:		data <= 32'h00000000;
		12'h7dc:		data <= 32'h0c000b23;
		12'h7dd:		data <= 32'h00000000;
		12'h7de:		data <= 32'h401a6000;
		12'h7df:		data <= 32'h375a0004;
		12'h7e0:		data <= 32'h409a6000;
		12'h7e1:		data <= 32'h8fa80048;
		12'h7e2:		data <= 32'h8fa9004c;
		12'h7e3:		data <= 32'h8fba0050;
		12'h7e4:		data <= 32'h01000011;
		12'h7e5:		data <= 32'h01200013;
		12'h7e6:		data <= 32'h8fa10000;
		12'h7e7:		data <= 32'h8fa20004;
		12'h7e8:		data <= 32'h8fa30008;
		12'h7e9:		data <= 32'h8fa4000c;
		12'h7ea:		data <= 32'h8fa50010;
		12'h7eb:		data <= 32'h8fa60014;
		12'h7ec:		data <= 32'h8fa70018;
		12'h7ed:		data <= 32'h8fa8001c;
		12'h7ee:		data <= 32'h8fa90020;
		12'h7ef:		data <= 32'h8faa0024;
		12'h7f0:		data <= 32'h8fab0028;
		12'h7f1:		data <= 32'h8fac002c;
		12'h7f2:		data <= 32'h8fad0030;
		12'h7f3:		data <= 32'h8fae0034;
		12'h7f4:		data <= 32'h8faf0038;
		12'h7f5:		data <= 32'h8fb8003c;
		12'h7f6:		data <= 32'h8fb90040;
		12'h7f7:		data <= 32'h8fbf0044;
		12'h7f8:		data <= 32'h27bd0054;
		12'h7f9:		data <= 32'h03400008;
		12'h7fa:		data <= 32'h42000010;
		12'h7fb:		data <= 32'h3c02f000;
		12'h7fc:		data <= 32'hac400000;
		12'h7fd:		data <= 32'h34440014;
		12'h7fe:		data <= 32'h34430010;
		12'h7ff:		data <= 32'h8c630000;
		12'h800:		data <= 32'h8c850000;
		12'h801:		data <= 32'h00003021;
		12'h802:		data <= 32'h34440020;
		12'h803:		data <= 32'h24a5ffff;
		12'h804:		data <= 32'h24c60001;
		12'h805:		data <= 32'h0066102b;
		12'h806:		data <= 32'hac800000;
		12'h807:		data <= 32'hac800004;
		12'h808:		data <= 32'hac85000c;
		12'h809:		data <= 32'h1040fffa;
		12'h80a:		data <= 32'h24840010;
		12'h80b:		data <= 32'h24030001;
		12'h80c:		data <= 32'h3c02f000;
		12'h80d:		data <= 32'hac430000;
		12'h80e:		data <= 32'h03e00008;
		12'h80f:		data <= 32'h00000000;
		12'h810:		data <= 32'h3c020100;
		12'h811:		data <= 32'h8c4326bc;
		12'h812:		data <= 32'h27bdffe0;
		12'h813:		data <= 32'h30630009;
		12'h814:		data <= 32'hafb10014;
		12'h815:		data <= 32'hafb00010;
		12'h816:		data <= 32'hafbf0018;
		12'h817:		data <= 32'h00a08821;
		12'h818:		data <= 32'h14600003;
		12'h819:		data <= 32'h00808021;
		12'h81a:		data <= 32'h0c00078e;
		12'h81b:		data <= 32'h00000000;
		12'h81c:		data <= 32'h0220f809;
		12'h81d:		data <= 32'h02002021;
		12'h81e:		data <= 32'h8fbf0018;
		12'h81f:		data <= 32'h8fb10014;
		12'h820:		data <= 32'h8fb00010;
		12'h821:		data <= 32'h08000a36;
		12'h822:		data <= 32'h27bd0020;
		12'h823:		data <= 32'h27bdffe8;
		12'h824:		data <= 32'hafbf0010;
		12'h825:		data <= 32'h0c000b2f;
		12'h826:		data <= 32'h00000000;
		12'h827:		data <= 32'h0c000b2f;
		12'h828:		data <= 32'h00000000;
		12'h829:		data <= 32'h08000825;
		12'h82a:		data <= 32'h00000000;
		12'h82b:		data <= 32'h27bdffe8;
		12'h82c:		data <= 32'h3c060100;
		12'h82d:		data <= 32'hafbf0014;
		12'h82e:		data <= 32'hafb00010;
		12'h82f:		data <= 32'h24c32698;
		12'h830:		data <= 32'h8c620024;
		12'h831:		data <= 32'h00000000;
		12'h832:		data <= 32'h10400006;
		12'h833:		data <= 32'h24020001;
		12'h834:		data <= 32'ha0620028;
		12'h835:		data <= 32'h8fbf0014;
		12'h836:		data <= 32'h8fb00010;
		12'h837:		data <= 32'h03e00008;
		12'h838:		data <= 32'h27bd0018;
		12'h839:		data <= 32'h8cc22698;
		12'h83a:		data <= 32'h00000000;
		12'h83b:		data <= 32'h14400018;
		12'h83c:		data <= 32'ha0600028;
		12'h83d:		data <= 32'h00003821;
		12'h83e:		data <= 32'h24c22698;
		12'h83f:		data <= 32'h8c50002c;
		12'h840:		data <= 32'h00000000;
		12'h841:		data <= 32'h10f0fff3;
		12'h842:		data <= 32'h00000000;
		12'h843:		data <= 32'h14e0001f;
		12'h844:		data <= 32'h3c020100;
		12'h845:		data <= 32'h3c020100;
		12'h846:		data <= 32'h244426c8;
		12'h847:		data <= 32'h16000015;
		12'h848:		data <= 32'h3c020100;
		12'h849:		data <= 32'h3c020100;
		12'h84a:		data <= 32'h244526c8;
		12'h84b:		data <= 32'h24c22698;
		12'h84c:		data <= 32'h0c0007a4;
		12'h84d:		data <= 32'hac47002c;
		12'h84e:		data <= 32'h1200ffe6;
		12'h84f:		data <= 32'h02002021;
		12'h850:		data <= 32'h8fbf0014;
		12'h851:		data <= 32'h8fb00010;
		12'h852:		data <= 32'h08000a7a;
		12'h853:		data <= 32'h27bd0018;
		12'h854:		data <= 32'h3c030100;
		12'h855:		data <= 32'h00021080;
		12'h856:		data <= 32'h24630078;
		12'h857:		data <= 32'h00431021;
		12'h858:		data <= 32'h8c44fffc;
		12'h859:		data <= 32'h00000000;
		12'h85a:		data <= 32'h8c870008;
		12'h85b:		data <= 32'h0800083f;
		12'h85c:		data <= 32'h24c22698;
		12'h85d:		data <= 32'h00101880;
		12'h85e:		data <= 32'h24420078;
		12'h85f:		data <= 32'h00621821;
		12'h860:		data <= 32'h8c65fffc;
		12'h861:		data <= 32'h0800084c;
		12'h862:		data <= 32'h24c22698;
		12'h863:		data <= 32'h00071880;
		12'h864:		data <= 32'h24420078;
		12'h865:		data <= 32'h00621821;
		12'h866:		data <= 32'h8c64fffc;
		12'h867:		data <= 32'h08000847;
		12'h868:		data <= 32'h00000000;
		12'h869:		data <= 32'h3c020100;
		12'h86a:		data <= 32'h00041880;
		12'h86b:		data <= 32'h24420078;
		12'h86c:		data <= 32'h00621821;
		12'h86d:		data <= 32'h00802821;
		12'h86e:		data <= 32'h8c64fffc;
		12'h86f:		data <= 32'h24020002;
		12'h870:		data <= 32'ha0820018;
		12'h871:		data <= 32'h3c040100;
		12'h872:		data <= 32'h080008b3;
		12'h873:		data <= 32'h24842698;
		12'h874:		data <= 32'h3c020100;
		12'h875:		data <= 32'h00041880;
		12'h876:		data <= 32'h24420078;
		12'h877:		data <= 32'h00621821;
		12'h878:		data <= 32'h00802821;
		12'h879:		data <= 32'h8c64fffc;
		12'h87a:		data <= 32'h24020004;
		12'h87b:		data <= 32'ha0820018;
		12'h87c:		data <= 32'h3c040100;
		12'h87d:		data <= 32'h080008de;
		12'h87e:		data <= 32'h24842698;
		12'h87f:		data <= 32'h3c020100;
		12'h880:		data <= 32'h27bdffe8;
		12'h881:		data <= 32'h00041880;
		12'h882:		data <= 32'h24420078;
		12'h883:		data <= 32'h00621821;
		12'h884:		data <= 32'hafbf0014;
		12'h885:		data <= 32'hafb00010;
		12'h886:		data <= 32'h8c70fffc;
		12'h887:		data <= 32'h00802821;
		12'h888:		data <= 32'h92020018;
		12'h889:		data <= 32'h3c040100;
		12'h88a:		data <= 32'h30420008;
		12'h88b:		data <= 32'h24842698;
		12'h88c:		data <= 32'h14400004;
		12'h88d:		data <= 32'h24030008;
		12'h88e:		data <= 32'h0c0008b3;
		12'h88f:		data <= 32'h00000000;
		12'h890:		data <= 32'h24030002;
		12'h891:		data <= 32'ha2030018;
		12'h892:		data <= 32'h8fbf0014;
		12'h893:		data <= 32'h8fb00010;
		12'h894:		data <= 32'h03e00008;
		12'h895:		data <= 32'h27bd0018;
		12'h896:		data <= 32'h30c60001;
		12'h897:		data <= 32'h10c00003;
		12'h898:		data <= 32'h00000000;
		12'h899:		data <= 32'h080008b3;
		12'h89a:		data <= 32'h00000000;
		12'h89b:		data <= 32'h0800089d;
		12'h89c:		data <= 32'h00000000;
		12'h89d:		data <= 32'h3c030100;
		12'h89e:		data <= 32'h24630078;
		12'h89f:		data <= 32'h00051080;
		12'h8a0:		data <= 32'h00803821;
		12'h8a1:		data <= 32'h00431021;
		12'h8a2:		data <= 32'h8c840000;
		12'h8a3:		data <= 32'h8c46fffc;
		12'h8a4:		data <= 32'h00041080;
		12'h8a5:		data <= 32'hacc70004;
		12'h8a6:		data <= 32'h14800004;
		12'h8a7:		data <= 32'h00431021;
		12'h8a8:		data <= 32'hacc50008;
		12'h8a9:		data <= 32'h03e00008;
		12'h8aa:		data <= 32'hace50000;
		12'h8ab:		data <= 32'h8c43fffc;
		12'h8ac:		data <= 32'h00000000;
		12'h8ad:		data <= 32'h8c620008;
		12'h8ae:		data <= 32'h00000000;
		12'h8af:		data <= 32'hacc20008;
		12'h8b0:		data <= 32'hac650008;
		12'h8b1:		data <= 32'h03e00008;
		12'h8b2:		data <= 32'hace50000;
		12'h8b3:		data <= 32'h3c030100;
		12'h8b4:		data <= 32'h24630078;
		12'h8b5:		data <= 32'h00051080;
		12'h8b6:		data <= 32'h00431021;
		12'h8b7:		data <= 32'h8c4afffc;
		12'h8b8:		data <= 32'h8c890000;
		12'h8b9:		data <= 32'h00000000;
		12'h8ba:		data <= 32'h15200004;
		12'h8bb:		data <= 32'had440004;
		12'h8bc:		data <= 32'had450008;
		12'h8bd:		data <= 32'h03e00008;
		12'h8be:		data <= 32'hac850000;
		12'h8bf:		data <= 32'h00091080;
		12'h8c0:		data <= 32'h00431021;
		12'h8c1:		data <= 32'h8c48fffc;
		12'h8c2:		data <= 32'h00606021;
		12'h8c3:		data <= 32'h8d070008;
		12'h8c4:		data <= 32'h914b0019;
		12'h8c5:		data <= 32'h00071080;
		12'h8c6:		data <= 32'h00431021;
		12'h8c7:		data <= 32'h8c43fffc;
		12'h8c8:		data <= 32'h080008cc;
		12'h8c9:		data <= 32'h00000000;
		12'h8ca:		data <= 32'h00c03821;
		12'h8cb:		data <= 32'h00401821;
		12'h8cc:		data <= 32'h90620019;
		12'h8cd:		data <= 32'h00000000;
		12'h8ce:		data <= 32'h0162102a;
		12'h8cf:		data <= 32'h1440000b;
		12'h8d0:		data <= 32'h00000000;
		12'h8d1:		data <= 32'h8c660008;
		12'h8d2:		data <= 32'h00000000;
		12'h8d3:		data <= 32'h00061080;
		12'h8d4:		data <= 32'h004c1021;
		12'h8d5:		data <= 32'h8c42fffc;
		12'h8d6:		data <= 32'h14e9fff3;
		12'h8d7:		data <= 32'h00604021;
		12'h8d8:		data <= 32'hac850000;
		12'h8d9:		data <= 32'h00604021;
		12'h8da:		data <= 32'h00c03821;
		12'h8db:		data <= 32'had050008;
		12'h8dc:		data <= 32'h03e00008;
		12'h8dd:		data <= 32'had470008;
		12'h8de:		data <= 32'h3c030100;
		12'h8df:		data <= 32'h24630078;
		12'h8e0:		data <= 32'h00051080;
		12'h8e1:		data <= 32'h00431021;
		12'h8e2:		data <= 32'h8c4afffc;
		12'h8e3:		data <= 32'h00000000;
		12'h8e4:		data <= 32'h8d490008;
		12'h8e5:		data <= 32'h00000000;
		12'h8e6:		data <= 32'h10a90020;
		12'h8e7:		data <= 32'h00000000;
		12'h8e8:		data <= 32'h8c880000;
		12'h8e9:		data <= 32'h00000000;
		12'h8ea:		data <= 32'h00081080;
		12'h8eb:		data <= 32'h00431021;
		12'h8ec:		data <= 32'h8c46fffc;
		12'h8ed:		data <= 32'h00000000;
		12'h8ee:		data <= 32'h8cc70008;
		12'h8ef:		data <= 32'h00000000;
		12'h8f0:		data <= 32'h14a70005;
		12'h8f1:		data <= 32'h00071080;
		12'h8f2:		data <= 32'h080008fe;
		12'h8f3:		data <= 32'hacc90008;
		12'h8f4:		data <= 32'h00403821;
		12'h8f5:		data <= 32'h00071080;
		12'h8f6:		data <= 32'h00431021;
		12'h8f7:		data <= 32'h8c46fffc;
		12'h8f8:		data <= 32'h00000000;
		12'h8f9:		data <= 32'h8cc20008;
		12'h8fa:		data <= 32'h00000000;
		12'h8fb:		data <= 32'h1445fff8;
		12'h8fc:		data <= 32'h00e04021;
		12'h8fd:		data <= 32'hacc90008;
		12'h8fe:		data <= 32'h8c820000;
		12'h8ff:		data <= 32'h00000000;
		12'h900:		data <= 32'h10a20003;
		12'h901:		data <= 32'h00000000;
		12'h902:		data <= 32'h03e00008;
		12'h903:		data <= 32'had400004;
		12'h904:		data <= 32'hac880000;
		12'h905:		data <= 32'h03e00008;
		12'h906:		data <= 32'had400004;
		12'h907:		data <= 32'hac800000;
		12'h908:		data <= 32'h03e00008;
		12'h909:		data <= 32'had400004;
		12'h90a:		data <= 32'h8c830000;
		12'h90b:		data <= 32'h3c020100;
		12'h90c:		data <= 32'h24450078;
		12'h90d:		data <= 32'h00031080;
		12'h90e:		data <= 32'h00003021;
		12'h90f:		data <= 32'h1060000d;
		12'h910:		data <= 32'h00451021;
		12'h911:		data <= 32'h8c47fffc;
		12'h912:		data <= 32'h00000000;
		12'h913:		data <= 32'h8ce60008;
		12'h914:		data <= 32'h00000000;
		12'h915:		data <= 32'h00061080;
		12'h916:		data <= 32'h00451021;
		12'h917:		data <= 32'h8c45fffc;
		12'h918:		data <= 32'h10660006;
		12'h919:		data <= 32'h00000000;
		12'h91a:		data <= 32'h8ca20008;
		12'h91b:		data <= 32'haca00004;
		12'h91c:		data <= 32'hace20008;
		12'h91d:		data <= 32'h03e00008;
		12'h91e:		data <= 32'h00c01021;
		12'h91f:		data <= 32'hac800000;
		12'h920:		data <= 32'h0800091d;
		12'h921:		data <= 32'haca00004;
		12'h922:		data <= 32'h8c820000;
		12'h923:		data <= 32'h90880005;
		12'h924:		data <= 32'h90830004;
		12'h925:		data <= 32'h01021021;
		12'h926:		data <= 32'hac820000;
		12'h927:		data <= 32'h8ca60004;
		12'h928:		data <= 32'h00000000;
		12'h929:		data <= 32'h0066102b;
		12'h92a:		data <= 32'h1040000b;
		12'h92b:		data <= 32'h00000000;
		12'h92c:		data <= 32'h8ca20000;
		12'h92d:		data <= 32'h24630001;
		12'h92e:		data <= 32'h24450001;
		12'h92f:		data <= 32'h0066102b;
		12'h930:		data <= 32'h1440000a;
		12'h931:		data <= 32'h00003821;
		12'h932:		data <= 32'h01001021;
		12'h933:		data <= 32'ha0850005;
		12'h934:		data <= 32'h03e00008;
		12'h935:		data <= 32'ha0870004;
		12'h936:		data <= 32'h24630001;
		12'h937:		data <= 32'h0066102b;
		12'h938:		data <= 32'h8ca50000;
		12'h939:		data <= 32'h1040fff8;
		12'h93a:		data <= 32'h00003821;
		12'h93b:		data <= 32'h306700ff;
		12'h93c:		data <= 32'h01001021;
		12'h93d:		data <= 32'ha0850005;
		12'h93e:		data <= 32'h03e00008;
		12'h93f:		data <= 32'ha0870004;
		12'h940:		data <= 32'h27bdffd8;
		12'h941:		data <= 32'hafb40020;
		12'h942:		data <= 32'hafb20018;
		12'h943:		data <= 32'hafbf0024;
		12'h944:		data <= 32'hafb3001c;
		12'h945:		data <= 32'hafb10014;
		12'h946:		data <= 32'hafb00010;
		12'h947:		data <= 32'h8c910000;
		12'h948:		data <= 32'h0080a021;
		12'h949:		data <= 32'h1220000e;
		12'h94a:		data <= 32'h00a09021;
		12'h94b:		data <= 32'h3c130100;
		12'h94c:		data <= 32'h26630078;
		12'h94d:		data <= 32'h00111080;
		12'h94e:		data <= 32'h00431021;
		12'h94f:		data <= 32'h8c50fffc;
		12'h950:		data <= 32'h00000000;
		12'h951:		data <= 32'h8e030014;
		12'h952:		data <= 32'h00000000;
		12'h953:		data <= 32'h00a3102b;
		12'h954:		data <= 32'h1040000b;
		12'h955:		data <= 32'h00721023;
		12'h956:		data <= 32'hae020014;
		12'h957:		data <= 32'hae910000;
		12'h958:		data <= 32'h8fbf0024;
		12'h959:		data <= 32'h8fb40020;
		12'h95a:		data <= 32'h8fb3001c;
		12'h95b:		data <= 32'h8fb20018;
		12'h95c:		data <= 32'h8fb10014;
		12'h95d:		data <= 32'h8fb00010;
		12'h95e:		data <= 32'h03e00008;
		12'h95f:		data <= 32'h27bd0028;
		12'h960:		data <= 32'h2402ffce;
		12'h961:		data <= 32'ha2020024;
		12'h962:		data <= 32'h02202021;
		12'h963:		data <= 32'h0c00087f;
		12'h964:		data <= 32'h02439023;
		12'h965:		data <= 32'h0c00082b;
		12'h966:		data <= 32'h00000000;
		12'h967:		data <= 32'h8e05000c;
		12'h968:		data <= 32'h8e060010;
		12'h969:		data <= 32'h24a2ffff;
		12'h96a:		data <= 32'h26640078;
		12'h96b:		data <= 32'h00021080;
		12'h96c:		data <= 32'h00061880;
		12'h96d:		data <= 32'h00441021;
		12'h96e:		data <= 32'h00641821;
		12'h96f:		data <= 32'h8c420000;
		12'h970:		data <= 32'h8c64fffc;
		12'h971:		data <= 32'h10b1000c;
		12'h972:		data <= 32'h00008821;
		12'h973:		data <= 32'h8c430014;
		12'h974:		data <= 32'hac460010;
		12'h975:		data <= 32'hae000010;
		12'h976:		data <= 32'h00408021;
		12'h977:		data <= 32'h0243102b;
		12'h978:		data <= 32'hac85000c;
		12'h979:		data <= 32'h1040ffe6;
		12'h97a:		data <= 32'h00a08821;
		12'h97b:		data <= 32'h00721023;
		12'h97c:		data <= 32'h08000957;
		12'h97d:		data <= 32'hae020014;
		12'h97e:		data <= 32'h08000957;
		12'h97f:		data <= 32'hae000010;
		12'h980:		data <= 32'h3c020100;
		12'h981:		data <= 32'h24470078;
		12'h982:		data <= 32'h00051880;
		12'h983:		data <= 32'h8c8a0000;
		12'h984:		data <= 32'h00671821;
		12'h985:		data <= 32'h8c6bfffc;
		12'h986:		data <= 32'h15400006;
		12'h987:		data <= 32'h00e07021;
		12'h988:		data <= 32'had65000c;
		12'h989:		data <= 32'had650010;
		12'h98a:		data <= 32'had660014;
		12'h98b:		data <= 32'h03e00008;
		12'h98c:		data <= 32'hac850000;
		12'h98d:		data <= 32'h000a1080;
		12'h98e:		data <= 32'h00471021;
		12'h98f:		data <= 32'h8c48fffc;
		12'h990:		data <= 32'h08000994;
		12'h991:		data <= 32'h01404821;
		12'h992:		data <= 32'h00604821;
		12'h993:		data <= 32'h00404021;
		12'h994:		data <= 32'h8d070014;
		12'h995:		data <= 32'h00000000;
		12'h996:		data <= 32'h00c7102b;
		12'h997:		data <= 32'h1440000f;
		12'h998:		data <= 32'h00000000;
		12'h999:		data <= 32'h8d03000c;
		12'h99a:		data <= 32'h00c73023;
		12'h99b:		data <= 32'h00031080;
		12'h99c:		data <= 32'h004e1021;
		12'h99d:		data <= 32'h01006821;
		12'h99e:		data <= 32'h8c42fffc;
		12'h99f:		data <= 32'h1543fff2;
		12'h9a0:		data <= 32'h01206021;
		12'h9a1:		data <= 32'had690010;
		12'h9a2:		data <= 32'had6a000c;
		12'h9a3:		data <= 32'hac450010;
		12'h9a4:		data <= 32'had660014;
		12'h9a5:		data <= 32'h03e00008;
		12'h9a6:		data <= 32'had05000c;
		12'h9a7:		data <= 32'h11490009;
		12'h9a8:		data <= 32'h00000000;
		12'h9a9:		data <= 32'h00e61023;
		12'h9aa:		data <= 32'had6c0010;
		12'h9ab:		data <= 32'had020014;
		12'h9ac:		data <= 32'had69000c;
		12'h9ad:		data <= 32'had050010;
		12'h9ae:		data <= 32'had660014;
		12'h9af:		data <= 32'h03e00008;
		12'h9b0:		data <= 32'hada5000c;
		12'h9b1:		data <= 32'hac850000;
		12'h9b2:		data <= 32'h8d0c0010;
		12'h9b3:		data <= 32'h00000000;
		12'h9b4:		data <= 32'h000c1080;
		12'h9b5:		data <= 32'h004e1021;
		12'h9b6:		data <= 32'h8c4dfffc;
		12'h9b7:		data <= 32'h080009aa;
		12'h9b8:		data <= 32'h00e61023;
		12'h9b9:		data <= 32'h3c030100;
		12'h9ba:		data <= 32'h24630078;
		12'h9bb:		data <= 32'h00051080;
		12'h9bc:		data <= 32'h00431021;
		12'h9bd:		data <= 32'h8c49fffc;
		12'h9be:		data <= 32'h00000000;
		12'h9bf:		data <= 32'h8d260010;
		12'h9c0:		data <= 32'h00000000;
		12'h9c1:		data <= 32'h10c00015;
		12'h9c2:		data <= 32'h00061080;
		12'h9c3:		data <= 32'h10a60015;
		12'h9c4:		data <= 32'h00431021;
		12'h9c5:		data <= 32'h8d28000c;
		12'h9c6:		data <= 32'h8c4bfffc;
		12'h9c7:		data <= 32'h8c8a0000;
		12'h9c8:		data <= 32'h00081080;
		12'h9c9:		data <= 32'h00431021;
		12'h9ca:		data <= 32'h8c47fffc;
		12'h9cb:		data <= 32'h110a0006;
		12'h9cc:		data <= 32'h00000000;
		12'h9cd:		data <= 32'h8ce20014;
		12'h9ce:		data <= 32'h8d230014;
		12'h9cf:		data <= 32'h00000000;
		12'h9d0:		data <= 32'h00431021;
		12'h9d1:		data <= 32'hace20014;
		12'h9d2:		data <= 32'h10aa0009;
		12'h9d3:		data <= 32'h00000000;
		12'h9d4:		data <= 32'had68000c;
		12'h9d5:		data <= 32'hace60010;
		12'h9d6:		data <= 32'had200010;
		12'h9d7:		data <= 32'h03e00008;
		12'h9d8:		data <= 32'h00000000;
		12'h9d9:		data <= 32'hac800000;
		12'h9da:		data <= 32'h03e00008;
		12'h9db:		data <= 32'had200010;
		12'h9dc:		data <= 32'hac880000;
		12'h9dd:		data <= 32'had68000c;
		12'h9de:		data <= 32'h080009d6;
		12'h9df:		data <= 32'hace60010;
		12'h9e0:		data <= 32'h27bdffe0;
		12'h9e1:		data <= 32'hafb10014;
		12'h9e2:		data <= 32'hafb00010;
		12'h9e3:		data <= 32'hafbf0018;
		12'h9e4:		data <= 32'h8c880000;
		12'h9e5:		data <= 32'h00808021;
		12'h9e6:		data <= 32'h1100001f;
		12'h9e7:		data <= 32'h00a08821;
		12'h9e8:		data <= 32'h01001821;
		12'h9e9:		data <= 32'h080009ed;
		12'h9ea:		data <= 32'hae080008;
		12'h9eb:		data <= 32'h10680018;
		12'h9ec:		data <= 32'hacc70008;
		12'h9ed:		data <= 32'h8c620000;
		12'h9ee:		data <= 32'h00603021;
		12'h9ef:		data <= 32'hae020004;
		12'h9f0:		data <= 32'h8c620008;
		12'h9f1:		data <= 32'h00602021;
		12'h9f2:		data <= 32'h8c630000;
		12'h9f3:		data <= 32'h02222823;
		12'h9f4:		data <= 32'h00513823;
		12'h9f5:		data <= 32'h0222102b;
		12'h9f6:		data <= 32'h1440fff4;
		12'h9f7:		data <= 32'hae030008;
		12'h9f8:		data <= 32'h8cc2000c;
		12'h9f9:		data <= 32'h00000000;
		12'h9fa:		data <= 32'h0040f809;
		12'h9fb:		data <= 32'h00000000;
		12'h9fc:		data <= 32'h8e030008;
		12'h9fd:		data <= 32'h00000000;
		12'h9fe:		data <= 32'h10600005;
		12'h9ff:		data <= 32'h00000000;
		12'ha00:		data <= 32'h8e080000;
		12'ha01:		data <= 32'h00000000;
		12'ha02:		data <= 32'h1468ffea;
		12'ha03:		data <= 32'h00000000;
		12'ha04:		data <= 32'hae000004;
		12'ha05:		data <= 32'hae000008;
		12'ha06:		data <= 32'h8fbf0018;
		12'ha07:		data <= 32'h8fb10014;
		12'ha08:		data <= 32'h8fb00010;
		12'ha09:		data <= 32'h03e00008;
		12'ha0a:		data <= 32'h27bd0020;
		12'ha0b:		data <= 32'h8c860000;
		12'ha0c:		data <= 32'h00000000;
		12'ha0d:		data <= 32'h14c00004;
		12'ha0e:		data <= 32'h24a3001f;
		12'ha0f:		data <= 32'h00001821;
		12'ha10:		data <= 32'h03e00008;
		12'ha11:		data <= 32'h00601021;
		12'ha12:		data <= 32'h8cc40004;
		12'ha13:		data <= 32'h2402ffe0;
		12'ha14:		data <= 32'h1080fffa;
		12'ha15:		data <= 32'h00624024;
		12'ha16:		data <= 32'h3405abcd;
		12'ha17:		data <= 32'h8cc70008;
		12'ha18:		data <= 32'h00861821;
		12'ha19:		data <= 32'h14e50003;
		12'ha1a:		data <= 32'h0088102b;
		12'ha1b:		data <= 32'h10400008;
		12'ha1c:		data <= 32'h00000000;
		12'ha1d:		data <= 32'h24660020;
		12'ha1e:		data <= 32'h8cc40004;
		12'ha1f:		data <= 32'h00000000;
		12'ha20:		data <= 32'h1480fff6;
		12'ha21:		data <= 32'h00001821;
		12'ha22:		data <= 32'h08000a10;
		12'ha23:		data <= 32'h00000000;
		12'ha24:		data <= 32'h00882823;
		12'ha25:		data <= 32'h2ca20041;
		12'ha26:		data <= 32'h1440000b;
		12'ha27:		data <= 32'h24c30020;
		12'ha28:		data <= 32'h00c81821;
		12'ha29:		data <= 32'h24620020;
		12'ha2a:		data <= 32'h24a5ffe0;
		12'ha2b:		data <= 32'h00c42021;
		12'ha2c:		data <= 32'hac660020;
		12'ha2d:		data <= 32'hac450004;
		12'ha2e:		data <= 32'hac820020;
		12'ha2f:		data <= 32'hac470008;
		12'ha30:		data <= 32'hacc80004;
		12'ha31:		data <= 32'h24c30020;
		12'ha32:		data <= 32'h24021234;
		12'ha33:		data <= 32'hacc20008;
		12'ha34:		data <= 32'h03e00008;
		12'ha35:		data <= 32'h00601021;
		12'ha36:		data <= 32'h27bdffe0;
		12'ha37:		data <= 32'h3c020100;
		12'ha38:		data <= 32'hafbf0018;
		12'ha39:		data <= 32'hafb00010;
		12'ha3a:		data <= 32'hafb10014;
		12'ha3b:		data <= 32'h8c5126c4;
		12'ha3c:		data <= 32'h0c000786;
		12'ha3d:		data <= 32'h00000000;
		12'ha3e:		data <= 32'h0c000b50;
		12'ha3f:		data <= 32'h02202021;
		12'ha40:		data <= 32'h3c020100;
		12'ha41:		data <= 32'h00111880;
		12'ha42:		data <= 32'h24420078;
		12'ha43:		data <= 32'h00621821;
		12'ha44:		data <= 32'h8c70fffc;
		12'ha45:		data <= 32'h00000000;
		12'ha46:		data <= 32'h8e040020;
		12'ha47:		data <= 32'h00000000;
		12'ha48:		data <= 32'h14800011;
		12'ha49:		data <= 32'h00000000;
		12'ha4a:		data <= 32'h9202001d;
		12'ha4b:		data <= 32'h00000000;
		12'ha4c:		data <= 32'h1440001b;
		12'ha4d:		data <= 32'h2442ffff;
		12'ha4e:		data <= 32'h0c00082b;
		12'ha4f:		data <= 32'ha2000018;
		12'ha50:		data <= 32'h8e070040;
		12'ha51:		data <= 32'h8e040034;
		12'ha52:		data <= 32'h8e050038;
		12'ha53:		data <= 32'h3c060000;
		12'ha54:		data <= 32'h8fbf0018;
		12'ha55:		data <= 32'h8fb10014;
		12'ha56:		data <= 32'h8fb00010;
		12'ha57:		data <= 32'h24c62040;
		12'ha58:		data <= 32'h08000b31;
		12'ha59:		data <= 32'h27bd0020;
		12'ha5a:		data <= 32'h0c000abd;
		12'ha5b:		data <= 32'h02202821;
		12'ha5c:		data <= 32'h8e040020;
		12'ha5d:		data <= 32'h00000000;
		12'ha5e:		data <= 32'h1080ffeb;
		12'ha5f:		data <= 32'h00000000;
		12'ha60:		data <= 32'h0c000abd;
		12'ha61:		data <= 32'h02202821;
		12'ha62:		data <= 32'h8e040020;
		12'ha63:		data <= 32'h00000000;
		12'ha64:		data <= 32'h1480fff5;
		12'ha65:		data <= 32'h00000000;
		12'ha66:		data <= 32'h08000a4a;
		12'ha67:		data <= 32'h00000000;
		12'ha68:		data <= 32'h9203003c;
		12'ha69:		data <= 32'h02202021;
		12'ha6a:		data <= 32'ha202001d;
		12'ha6b:		data <= 32'ha203001a;
		12'ha6c:		data <= 32'h0c000869;
		12'ha6d:		data <= 32'ha2030019;
		12'ha6e:		data <= 32'h0c00082b;
		12'ha6f:		data <= 32'h00000000;
		12'ha70:		data <= 32'h8e070040;
		12'ha71:		data <= 32'h8e040034;
		12'ha72:		data <= 32'h8e050038;
		12'ha73:		data <= 32'h3c060000;
		12'ha74:		data <= 32'h8fbf0018;
		12'ha75:		data <= 32'h8fb10014;
		12'ha76:		data <= 32'h8fb00010;
		12'ha77:		data <= 32'h24c62040;
		12'ha78:		data <= 32'h08000b31;
		12'ha79:		data <= 32'h27bd0020;
		12'ha7a:		data <= 32'h3c020100;
		12'ha7b:		data <= 32'h27bdffd8;
		12'ha7c:		data <= 32'h24420078;
		12'ha7d:		data <= 32'h00042080;
		12'ha7e:		data <= 32'hafbf0024;
		12'ha7f:		data <= 32'hafb40020;
		12'ha80:		data <= 32'hafb3001c;
		12'ha81:		data <= 32'hafb20018;
		12'ha82:		data <= 32'hafb10014;
		12'ha83:		data <= 32'hafb00010;
		12'ha84:		data <= 32'h00822021;
		12'ha85:		data <= 32'h8c90fffc;
		12'ha86:		data <= 32'h24020001;
		12'ha87:		data <= 32'h9203002c;
		12'ha88:		data <= 32'h00000000;
		12'ha89:		data <= 32'h10620009;
		12'ha8a:		data <= 32'h00000000;
		12'ha8b:		data <= 32'h8fbf0024;
		12'ha8c:		data <= 32'h8fb40020;
		12'ha8d:		data <= 32'h8fb3001c;
		12'ha8e:		data <= 32'h8fb20018;
		12'ha8f:		data <= 32'h8fb10014;
		12'ha90:		data <= 32'h8fb00010;
		12'ha91:		data <= 32'h03e00008;
		12'ha92:		data <= 32'h27bd0028;
		12'ha93:		data <= 32'h8e110030;
		12'ha94:		data <= 32'h00000000;
		12'ha95:		data <= 32'h1220fff5;
		12'ha96:		data <= 32'h3c020100;
		12'ha97:		data <= 32'h8e130034;
		12'ha98:		data <= 32'h08000aa2;
		12'ha99:		data <= 32'h24542698;
		12'ha9a:		data <= 32'h0240f809;
		12'ha9b:		data <= 32'h02602821;
		12'ha9c:		data <= 32'h0c000786;
		12'ha9d:		data <= 32'h00000000;
		12'ha9e:		data <= 32'h8e110030;
		12'ha9f:		data <= 32'h00000000;
		12'haa0:		data <= 32'h12200013;
		12'haa1:		data <= 32'h24020001;
		12'haa2:		data <= 32'ha200002c;
		12'haa3:		data <= 32'h8e820024;
		12'haa4:		data <= 32'hae000030;
		12'haa5:		data <= 32'h30420009;
		12'haa6:		data <= 32'h8e120044;
		12'haa7:		data <= 32'h1440fff2;
		12'haa8:		data <= 32'h3224ffff;
		12'haa9:		data <= 32'h0c00078e;
		12'haaa:		data <= 32'h00000000;
		12'haab:		data <= 32'h3224ffff;
		12'haac:		data <= 32'h0240f809;
		12'haad:		data <= 32'h02602821;
		12'haae:		data <= 32'h0c000786;
		12'haaf:		data <= 32'h00000000;
		12'hab0:		data <= 32'h8e110030;
		12'hab1:		data <= 32'h00000000;
		12'hab2:		data <= 32'h1620ffef;
		12'hab3:		data <= 32'h24020001;
		12'hab4:		data <= 32'ha202002c;
		12'hab5:		data <= 32'h8fbf0024;
		12'hab6:		data <= 32'h8fb40020;
		12'hab7:		data <= 32'h8fb3001c;
		12'hab8:		data <= 32'h8fb20018;
		12'hab9:		data <= 32'h8fb10014;
		12'haba:		data <= 32'h8fb00010;
		12'habb:		data <= 32'h03e00008;
		12'habc:		data <= 32'h27bd0028;
		12'habd:		data <= 32'h3c030100;
		12'habe:		data <= 32'h27bdffe0;
		12'habf:		data <= 32'h2469027c;
		12'hac0:		data <= 32'h00041080;
		12'hac1:		data <= 32'hafb20018;
		12'hac2:		data <= 32'hafb00010;
		12'hac3:		data <= 32'hafbf001c;
		12'hac4:		data <= 32'hafb10014;
		12'hac5:		data <= 32'h00491021;
		12'hac6:		data <= 32'h8c48fffc;
		12'hac7:		data <= 32'h3c120100;
		12'hac8:		data <= 32'h8d060008;
		12'hac9:		data <= 32'h00052880;
		12'haca:		data <= 32'h26430078;
		12'hacb:		data <= 32'h00061080;
		12'hacc:		data <= 32'h00a32821;
		12'hacd:		data <= 32'h00808021;
		12'hace:		data <= 32'had000004;
		12'hacf:		data <= 32'h8ca7fffc;
		12'had0:		data <= 32'h1086002c;
		12'had1:		data <= 32'h00491021;
		12'had2:		data <= 32'h8c45fffc;
		12'had3:		data <= 32'h00000000;
		12'had4:		data <= 32'h8ca4000c;
		12'had5:		data <= 32'h00000000;
		12'had6:		data <= 32'h00041080;
		12'had7:		data <= 32'h00491021;
		12'had8:		data <= 32'h8c43fffc;
		12'had9:		data <= 32'h00000000;
		12'hada:		data <= 32'hac660008;
		12'hadb:		data <= 32'h8ce20020;
		12'hadc:		data <= 32'h00000000;
		12'hadd:		data <= 32'h12020021;
		12'hade:		data <= 32'h00000000;
		12'hadf:		data <= 32'h0c00090a;
		12'hae0:		data <= 32'h01002021;
		12'hae1:		data <= 32'h00408821;
		12'hae2:		data <= 32'h26430078;
		12'hae3:		data <= 32'h00021080;
		12'hae4:		data <= 32'h00431021;
		12'hae5:		data <= 32'h02002021;
		12'hae6:		data <= 32'h16200007;
		12'hae7:		data <= 32'h02202821;
		12'hae8:		data <= 32'h8fbf001c;
		12'hae9:		data <= 32'h8fb20018;
		12'haea:		data <= 32'h8fb10014;
		12'haeb:		data <= 32'h8fb00010;
		12'haec:		data <= 32'h03e00008;
		12'haed:		data <= 32'h27bd0020;
		12'haee:		data <= 32'h8c50fffc;
		12'haef:		data <= 32'h0c000b5b;
		12'haf0:		data <= 32'h00000000;
		12'haf1:		data <= 32'h02202021;
		12'haf2:		data <= 32'h0c00087f;
		12'haf3:		data <= 32'ha2000024;
		12'haf4:		data <= 32'h3c040100;
		12'haf5:		data <= 32'h02202821;
		12'haf6:		data <= 32'h8fbf001c;
		12'haf7:		data <= 32'h8fb20018;
		12'haf8:		data <= 32'h8fb10014;
		12'haf9:		data <= 32'h8fb00010;
		12'hafa:		data <= 32'h248426a4;
		12'hafb:		data <= 32'h080009b9;
		12'hafc:		data <= 32'h27bd0020;
		12'hafd:		data <= 32'h08000adf;
		12'hafe:		data <= 32'hace00020;
		12'haff:		data <= 32'h08000adf;
		12'hb00:		data <= 32'hace60020;
		12'hb01:		data <= 32'h3c030100;
		12'hb02:		data <= 32'h24632698;
		12'hb03:		data <= 32'h8c620024;
		12'hb04:		data <= 32'h00000000;
		12'hb05:		data <= 32'h34420004;
		12'hb06:		data <= 32'h03e00008;
		12'hb07:		data <= 32'hac620024;
		12'hb08:		data <= 32'h3c030100;
		12'hb09:		data <= 32'h27bdffe0;
		12'hb0a:		data <= 32'h00041080;
		12'hb0b:		data <= 32'h24630244;
		12'hb0c:		data <= 32'hafb10014;
		12'hb0d:		data <= 32'hafb00010;
		12'hb0e:		data <= 32'hafbf0018;
		12'hb0f:		data <= 32'h00438021;
		12'hb10:		data <= 32'h00808821;
		12'hb11:		data <= 32'h8e040000;
		12'hb12:		data <= 32'h00000000;
		12'hb13:		data <= 32'h1080000a;
		12'hb14:		data <= 32'h02202021;
		12'hb15:		data <= 32'h0c00078e;
		12'hb16:		data <= 32'h00000000;
		12'hb17:		data <= 32'h8e020000;
		12'hb18:		data <= 32'h00000000;
		12'hb19:		data <= 32'h0040f809;
		12'hb1a:		data <= 32'h00000000;
		12'hb1b:		data <= 32'h0c000786;
		12'hb1c:		data <= 32'h00000000;
		12'hb1d:		data <= 32'h02202021;
		12'hb1e:		data <= 32'h8fbf0018;
		12'hb1f:		data <= 32'h8fb10014;
		12'hb20:		data <= 32'h8fb00010;
		12'hb21:		data <= 32'h08000b33;
		12'hb22:		data <= 32'h27bd0020;
		12'hb23:		data <= 32'h3c020100;
		12'hb24:		data <= 32'h24422698;
		12'hb25:		data <= 32'h8c430024;
		12'hb26:		data <= 32'h2404fffb;
		12'hb27:		data <= 32'h90450028;
		12'hb28:		data <= 32'h00641824;
		12'hb29:		data <= 32'h14a00003;
		12'hb2a:		data <= 32'hac430024;
		12'hb2b:		data <= 32'h03e00008;
		12'hb2c:		data <= 32'h00000000;
		12'hb2d:		data <= 32'h0800082b;
		12'hb2e:		data <= 32'h00000000;
		12'hb2f:		data <= 32'h1000ffff;
		12'hb30:		data <= 32'h00000000;
		12'hb31:		data <= 32'h00c00008;
		12'hb32:		data <= 32'h00e0e821;
		12'hb33:		data <= 32'h27bdffd8;
		12'hb34:		data <= 32'hafb00010;
		12'hb35:		data <= 32'h3c10f000;
		12'hb36:		data <= 32'hafbf0020;
		12'hb37:		data <= 32'hafb20018;
		12'hb38:		data <= 32'hafb10014;
		12'hb39:		data <= 32'hafb3001c;
		12'hb3a:		data <= 32'h36020008;
		12'hb3b:		data <= 32'hae000000;
		12'hb3c:		data <= 32'h8c440000;
		12'hb3d:		data <= 32'h36110004;
		12'hb3e:		data <= 32'h3602000c;
		12'hb3f:		data <= 32'h8e330000;
		12'hb40:		data <= 32'h8c430000;
		12'hb41:		data <= 32'h24120001;
		12'hb42:		data <= 32'hae230000;
		12'hb43:		data <= 32'hae120000;
		12'hb44:		data <= 32'h0c000b7a;
		12'hb45:		data <= 32'h00000000;
		12'hb46:		data <= 32'hae000000;
		12'hb47:		data <= 32'hae330000;
		12'hb48:		data <= 32'hae120000;
		12'hb49:		data <= 32'h8fbf0020;
		12'hb4a:		data <= 32'h8fb3001c;
		12'hb4b:		data <= 32'h8fb20018;
		12'hb4c:		data <= 32'h8fb10014;
		12'hb4d:		data <= 32'h8fb00010;
		12'hb4e:		data <= 32'h03e00008;
		12'hb4f:		data <= 32'h27bd0028;
		12'hb50:		data <= 32'h3c020100;
		12'hb51:		data <= 32'h00041880;
		12'hb52:		data <= 32'h24420078;
		12'hb53:		data <= 32'h00621821;
		12'hb54:		data <= 32'h00802821;
		12'hb55:		data <= 32'h8c64fffc;
		12'hb56:		data <= 32'h00000000;
		12'hb57:		data <= 32'ha0800018;
		12'hb58:		data <= 32'h3c040100;
		12'hb59:		data <= 32'h080008de;
		12'hb5a:		data <= 32'h24842698;
		12'hb5b:		data <= 32'h3c020100;
		12'hb5c:		data <= 32'h2447027c;
		12'hb5d:		data <= 32'h00804021;
		12'hb5e:		data <= 32'h3c020100;
		12'hb5f:		data <= 32'h00042080;
		12'hb60:		data <= 32'h00051880;
		12'hb61:		data <= 32'h24420078;
		12'hb62:		data <= 32'h00872021;
		12'hb63:		data <= 32'h00621821;
		12'hb64:		data <= 32'h8c86fffc;
		12'hb65:		data <= 32'h8c63fffc;
		12'hb66:		data <= 32'hacc50004;
		12'hb67:		data <= 32'h8c650020;
		12'hb68:		data <= 32'h00000000;
		12'hb69:		data <= 32'h00051080;
		12'hb6a:		data <= 32'h14a00004;
		12'hb6b:		data <= 32'h00471021;
		12'hb6c:		data <= 32'hac680020;
		12'hb6d:		data <= 32'h03e00008;
		12'hb6e:		data <= 32'hacc80008;
		12'hb6f:		data <= 32'h8c43fffc;
		12'hb70:		data <= 32'h00000000;
		12'hb71:		data <= 32'h8c64000c;
		12'hb72:		data <= 32'hac68000c;
		12'hb73:		data <= 32'h00041080;
		12'hb74:		data <= 32'h00471021;
		12'hb75:		data <= 32'h8c43fffc;
		12'hb76:		data <= 32'hacc4000c;
		12'hb77:		data <= 32'hac680008;
		12'hb78:		data <= 32'h03e00008;
		12'hb79:		data <= 32'hacc50008;
		12'hb7a:		data <= 32'h3c020000;
		12'hb7b:		data <= 32'h8c432e6c;
		12'hb7c:		data <= 32'h3c020100;
		12'hb7d:		data <= 32'h00832023;
		12'hb7e:		data <= 32'h27bdffe8;
		12'hb7f:		data <= 32'h00042080;
		12'hb80:		data <= 32'h24421288;
		12'hb81:		data <= 32'hafbf0014;
		12'hb82:		data <= 32'hafb00010;
		12'hb83:		data <= 32'h00822021;
		12'hb84:		data <= 32'h8c900000;
		12'hb85:		data <= 32'h00000000;
		12'hb86:		data <= 32'h1200000e;
		12'hb87:		data <= 32'h00000000;
		12'hb88:		data <= 32'h0c00078e;
		12'hb89:		data <= 32'h00000000;
		12'hb8a:		data <= 32'h8e040004;
		12'hb8b:		data <= 32'h8e020008;
		12'hb8c:		data <= 32'h00000000;
		12'hb8d:		data <= 32'h0040f809;
		12'hb8e:		data <= 32'h00000000;
		12'hb8f:		data <= 32'h0c000786;
		12'hb90:		data <= 32'h00000000;
		12'hb91:		data <= 32'h8e100000;
		12'hb92:		data <= 32'h00000000;
		12'hb93:		data <= 32'h1600fff4;
		12'hb94:		data <= 32'h00000000;
		12'hb95:		data <= 32'h8fbf0014;
		12'hb96:		data <= 32'h8fb00010;
		12'hb97:		data <= 32'h03e00008;
		12'hb98:		data <= 32'h27bd0018;
		12'hb99:		data <= 32'h00000004;
		12'hb9a:		data <= 32'h000000ff;
		12'hb9b:		data <= 32'h00000000;
		12'hb9c:		data <= 32'h00000000;
		12'hb9d:		data <= 32'h00000001;
		12'hb9e:		data <= 32'h00000000;
		12'hb9f:		data <= 32'h00000001;
		12'hba0:		data <= 32'h00000002;
		12'hba1:		data <= 32'h0000007f;
		12'hba2:		data <= 32'h00000002;
		12'hba3:		data <= 32'h00000002;
		12'hba4:		data <= 32'h00000006;
		12'hba5:		data <= 32'h00000006;
		12'hba6:		data <= 32'h01001288;
		12'hba7:		data <= 32'h7468696e;
		12'hba8:		data <= 32'h6b696e67;
		12'hba9:		data <= 32'h00000000;
		12'hbaa:		data <= 32'h68756e67;
		12'hbab:		data <= 32'h72790000;
		12'hbac:		data <= 32'h65617469;
		12'hbad:		data <= 32'h6e670000;
		12'hbae:		data <= 32'h01000068;
		12'hbaf:		data <= 32'h01000058;
		12'hbb0:		data <= 32'h01000048;
		12'hbb1:		data <= 32'h01000038;
		12'hbb2:		data <= 32'h01000028;
		12'hbb3:		data <= 32'h01000018;
		12'hbb4:		data <= 32'h00000000;
		12'hbb5:		data <= 32'h00000001;
		12'hbb6:		data <= 32'h00000000;
		12'hbb7:		data <= 32'h00000001;
		12'hbb8:		data <= 32'h00000000;
		12'hbb9:		data <= 32'h00000001;
		12'hbba:		data <= 32'h00000000;
		12'hbbb:		data <= 32'h00000001;
		12'hbbc:		data <= 32'h00000000;
		12'hbbd:		data <= 32'h00000001;
		12'hbbe:		data <= 32'h00000000;
		12'hbbf:		data <= 32'h00000001;
		12'hbc0:		data <= 32'h00000000;
		12'hbc1:		data <= 32'h00000001;
		12'hbc2:		data <= 32'h00000000;
		12'hbc3:		data <= 32'h00000001;
		12'hbc4:		data <= 32'h00000000;
		12'hbc5:		data <= 32'h00000001;
		12'hbc6:		data <= 32'h00000000;
		12'hbc7:		data <= 32'h00000001;
		12'hbc8:		data <= 32'h00000000;
		12'hbc9:		data <= 32'h00000001;
		12'hbca:		data <= 32'h00000000;
		12'hbcb:		data <= 32'h00000001;
		12'hbcc:		data <= 32'h010001f8;
		12'hbcd:		data <= 32'h010001b0;
		12'hbce:		data <= 32'h01000168;
		12'hbcf:		data <= 32'h01000120;
		12'hbd0:		data <= 32'h010000d8;
		12'hbd1:		data <= 32'h01000090;
		12'hbd2:		data <= 32'h00000000;
		12'hbd3:		data <= 32'h00000000;
		12'hbd4:		data <= 32'h00000000;
		12'hbd5:		data <= 32'h00000000;
		12'hbd6:		data <= 32'h00000000;
		12'hbd7:		data <= 32'h00000000;
		12'hbd8:		data <= 32'h00000000;
		12'hbd9:		data <= 32'h00000000;
		12'hbda:		data <= 32'h00000000;
		12'hbdb:		data <= 32'h00000000;
		12'hbdc:		data <= 32'h00000000;
		12'hbdd:		data <= 32'h00000000;
		12'hbde:		data <= 32'h00000000;
		12'hbdf:		data <= 32'h00000005;
		12'hbe0:		data <= 32'h0000048c;
		12'hbe1:		data <= 32'h02000000;
		12'hbe2:		data <= 32'h01000688;
		12'hbe3:		data <= 32'h00000000;
		12'hbe4:		data <= 32'h00000000;
		12'hbe5:		data <= 32'h00000000;
		12'hbe6:		data <= 32'h00000000;
		12'hbe7:		data <= 32'h00000000;
		12'hbe8:		data <= 32'h00000000;
		12'hbe9:		data <= 32'h00000000;
		12'hbea:		data <= 32'h00000000;
		12'hbeb:		data <= 32'h00000000;
		12'hbec:		data <= 32'h00000000;
		12'hbed:		data <= 32'h00000000;
		12'hbee:		data <= 32'h00000000;
		12'hbef:		data <= 32'h00000000;
		12'hbf0:		data <= 32'h00000000;
		12'hbf1:		data <= 32'h00000004;
		12'hbf2:		data <= 32'h0000048c;
		12'hbf3:		data <= 32'h02000000;
		12'hbf4:		data <= 32'h01000888;
		12'hbf5:		data <= 32'h00000000;
		12'hbf6:		data <= 32'h00000000;
		12'hbf7:		data <= 32'h00000000;
		12'hbf8:		data <= 32'h00000000;
		12'hbf9:		data <= 32'h00000000;
		12'hbfa:		data <= 32'h00000000;
		12'hbfb:		data <= 32'h00000000;
		12'hbfc:		data <= 32'h00000000;
		12'hbfd:		data <= 32'h00000000;
		12'hbfe:		data <= 32'h00000000;
		12'hbff:		data <= 32'h00000000;
		12'hc00:		data <= 32'h00000000;
		12'hc01:		data <= 32'h00000000;
		12'hc02:		data <= 32'h00000000;
		12'hc03:		data <= 32'h00000003;
		12'hc04:		data <= 32'h0000048c;
		12'hc05:		data <= 32'h02000000;
		12'hc06:		data <= 32'h01000a88;
		12'hc07:		data <= 32'h00000000;
		12'hc08:		data <= 32'h00000000;
		12'hc09:		data <= 32'h00000000;
		12'hc0a:		data <= 32'h00000000;
		12'hc0b:		data <= 32'h00000000;
		12'hc0c:		data <= 32'h00000000;
		12'hc0d:		data <= 32'h00000000;
		12'hc0e:		data <= 32'h00000000;
		12'hc0f:		data <= 32'h00000000;
		12'hc10:		data <= 32'h00000000;
		12'hc11:		data <= 32'h00000000;
		12'hc12:		data <= 32'h00000000;
		12'hc13:		data <= 32'h00000000;
		12'hc14:		data <= 32'h00000000;
		12'hc15:		data <= 32'h00000002;
		12'hc16:		data <= 32'h0000048c;
		12'hc17:		data <= 32'h02000000;
		12'hc18:		data <= 32'h01000c88;
		12'hc19:		data <= 32'h00000000;
		12'hc1a:		data <= 32'h00000000;
		12'hc1b:		data <= 32'h00000000;
		12'hc1c:		data <= 32'h00000000;
		12'hc1d:		data <= 32'h00000000;
		12'hc1e:		data <= 32'h00000000;
		12'hc1f:		data <= 32'h00000000;
		12'hc20:		data <= 32'h00000000;
		12'hc21:		data <= 32'h00000000;
		12'hc22:		data <= 32'h00000000;
		12'hc23:		data <= 32'h00000000;
		12'hc24:		data <= 32'h00000000;
		12'hc25:		data <= 32'h00000000;
		12'hc26:		data <= 32'h00000000;
		12'hc27:		data <= 32'h00000001;
		12'hc28:		data <= 32'h0000048c;
		12'hc29:		data <= 32'h02000000;
		12'hc2a:		data <= 32'h01000e88;
		12'hc2b:		data <= 32'h00000000;
		12'hc2c:		data <= 32'h00000000;
		12'hc2d:		data <= 32'h00000000;
		12'hc2e:		data <= 32'h00000000;
		12'hc2f:		data <= 32'h00000000;
		12'hc30:		data <= 32'h00000000;
		12'hc31:		data <= 32'h00000000;
		12'hc32:		data <= 32'h00000000;
		12'hc33:		data <= 32'h00000000;
		12'hc34:		data <= 32'h00000000;
		12'hc35:		data <= 32'h00000000;
		12'hc36:		data <= 32'h00000000;
		12'hc37:		data <= 32'h00000000;
		12'hc38:		data <= 32'h00000000;
		12'hc39:		data <= 32'h00000001;
		12'hc3a:		data <= 32'h0000060c;
		12'hc3b:		data <= 32'h01000000;
		12'hc3c:		data <= 32'h01001088;
		12'hc3d:		data <= 32'h00000000;
		12'hc3e:		data <= 32'h00003039;
		12'hc3f:		data <= 32'h00000000;
		12'hc40:		data <= 32'h00000000;
		12'hc41:		data <= 32'h00000000;
		12'hc42:		data <= 32'h00000000;
		12'hc43:		data <= 32'h00000000;
		12'hc44:		data <= 32'h00000000;
		12'hc45:		data <= 32'h00000000;
		12'hc46:		data <= 32'h00000000;
		12'hc47:		data <= 32'h00000000;
		12'hc48:		data <= 32'h00000000;
		12'hc49:		data <= 32'h00000000;
		12'hc4a:		data <= 32'h00000000;
		12'hc4b:		data <= 32'h00000000;
		12'hc4c:		data <= 32'h00000000;
		12'hc4d:		data <= 32'h00000000;
		12'hc4e:		data <= 32'h00000000;
		12'hc4f:		data <= 32'h00000000;
		12'hc50:		data <= 32'h00000000;
		12'hc51:		data <= 32'h00000000;
		12'hc52:		data <= 32'h00000000;
		12'hc53:		data <= 32'h00000000;
		12'hc54:		data <= 32'h00000000;
		12'hc55:		data <= 32'h00000000;
		12'hc56:		data <= 32'h00000000;
		12'hc57:		data <= 32'h00000000;
		12'hc58:		data <= 32'h00000000;
		12'hc59:		data <= 32'h00000000;
		12'hc5a:		data <= 32'h00000000;
		12'hc5b:		data <= 32'h00000000;
		12'hc5c:		data <= 32'h00000000;
		12'hc5d:		data <= 32'h00000000;
		12'hc5e:		data <= 32'h00000000;
		12'hc5f:		data <= 32'h00000000;
		12'hc60:		data <= 32'h00000000;
		12'hc61:		data <= 32'h00000000;
		12'hc62:		data <= 32'h00000000;
		12'hc63:		data <= 32'h00000000;
		12'hc64:		data <= 32'h00000000;
		12'hc65:		data <= 32'h00000000;
		12'hc66:		data <= 32'h00000000;
		12'hc67:		data <= 32'h00000000;
		12'hc68:		data <= 32'h00000000;
		12'hc69:		data <= 32'h00000000;
		12'hc6a:		data <= 32'h00000000;
		12'hc6b:		data <= 32'h00000000;
		12'hc6c:		data <= 32'h00000000;
		12'hc6d:		data <= 32'h00000000;
		12'hc6e:		data <= 32'h00000000;
		12'hc6f:		data <= 32'h00000000;
		12'hc70:		data <= 32'h00000000;
		12'hc71:		data <= 32'h00000000;
		12'hc72:		data <= 32'h00000000;
		12'hc73:		data <= 32'h00000000;
		12'hc74:		data <= 32'h00000000;
		12'hc75:		data <= 32'h00000000;
		12'hc76:		data <= 32'h00000000;
		12'hc77:		data <= 32'h00000000;
		12'hc78:		data <= 32'h00000000;
		12'hc79:		data <= 32'h00000000;
		12'hc7a:		data <= 32'h00000000;
		12'hc7b:		data <= 32'h00000000;
		12'hc7c:		data <= 32'h00000000;
		12'hc7d:		data <= 32'h00000000;
		12'hc7e:		data <= 32'h00000000;
		12'hc7f:		data <= 32'h00000000;
		12'hc80:		data <= 32'h00000000;
		12'hc81:		data <= 32'h00000000;
		12'hc82:		data <= 32'h00000000;
		12'hc83:		data <= 32'h00000000;
		12'hc84:		data <= 32'h00000000;
		12'hc85:		data <= 32'h00000000;
		12'hc86:		data <= 32'h00000000;
		12'hc87:		data <= 32'h00000000;
		12'hc88:		data <= 32'h00000000;
		12'hc89:		data <= 32'h00000000;
		12'hc8a:		data <= 32'h00000000;
		12'hc8b:		data <= 32'h00000000;
		12'hc8c:		data <= 32'h00000000;
		12'hc8d:		data <= 32'h00000000;
		12'hc8e:		data <= 32'h00000000;
		12'hc8f:		data <= 32'h00000000;
		12'hc90:		data <= 32'h00000000;
		12'hc91:		data <= 32'h00000000;
		12'hc92:		data <= 32'h00000000;
		12'hc93:		data <= 32'h00000000;
		12'hc94:		data <= 32'h00000000;
		12'hc95:		data <= 32'h00000000;
		12'hc96:		data <= 32'h00000000;
		12'hc97:		data <= 32'h00000000;
		12'hc98:		data <= 32'h00000000;
		12'hc99:		data <= 32'h00000000;
		12'hc9a:		data <= 32'h00000000;
		12'hc9b:		data <= 32'h00000000;
		12'hc9c:		data <= 32'h00000000;
		12'hc9d:		data <= 32'h00000000;
		12'hc9e:		data <= 32'h00000000;
		12'hc9f:		data <= 32'h00000000;
		12'hca0:		data <= 32'h00000000;
		12'hca1:		data <= 32'h00000000;
		12'hca2:		data <= 32'h00000000;
		12'hca3:		data <= 32'h00000000;
		12'hca4:		data <= 32'h00000000;
		12'hca5:		data <= 32'h00000000;
		12'hca6:		data <= 32'h00000000;
		12'hca7:		data <= 32'h00000000;
		12'hca8:		data <= 32'h00000000;
		12'hca9:		data <= 32'h00000000;
		12'hcaa:		data <= 32'h00000000;
		12'hcab:		data <= 32'h00000000;
		12'hcac:		data <= 32'h00000000;
		12'hcad:		data <= 32'h00000000;
		12'hcae:		data <= 32'h00000000;
		12'hcaf:		data <= 32'h00000000;
		12'hcb0:		data <= 32'h00000000;
		12'hcb1:		data <= 32'h00000000;
		12'hcb2:		data <= 32'h00000000;
		12'hcb3:		data <= 32'h00000000;
		12'hcb4:		data <= 32'h00000000;
		12'hcb5:		data <= 32'h00000000;
		12'hcb6:		data <= 32'h00000000;
		12'hcb7:		data <= 32'h00000000;
		12'hcb8:		data <= 32'h00000000;
		12'hcb9:		data <= 32'h00000000;
		12'hcba:		data <= 32'h00000000;
		12'hcbb:		data <= 32'h00000000;
		12'hcbc:		data <= 32'h00000000;
		12'hcbd:		data <= 32'h00000000;
		12'hcbe:		data <= 32'h00000000;
		12'hcbf:		data <= 32'h00000000;
		12'hcc0:		data <= 32'h00000000;
		12'hcc1:		data <= 32'h00000000;
		12'hcc2:		data <= 32'h00000000;
		12'hcc3:		data <= 32'h00000000;
		12'hcc4:		data <= 32'h00000000;
		12'hcc5:		data <= 32'h00000000;
		12'hcc6:		data <= 32'h00000000;
		12'hcc7:		data <= 32'h00000000;
		12'hcc8:		data <= 32'h00000000;
		12'hcc9:		data <= 32'h00000000;
		12'hcca:		data <= 32'h00000000;
		12'hccb:		data <= 32'h00000000;
		12'hccc:		data <= 32'h00000000;
		12'hccd:		data <= 32'h00000000;
		12'hcce:		data <= 32'h00000000;
		12'hccf:		data <= 32'h00000000;
		12'hcd0:		data <= 32'h00000000;
		12'hcd1:		data <= 32'h00000000;
		12'hcd2:		data <= 32'h00000000;
		12'hcd3:		data <= 32'h00000000;
		12'hcd4:		data <= 32'h00000000;
		12'hcd5:		data <= 32'h00000000;
		12'hcd6:		data <= 32'h00000000;
		12'hcd7:		data <= 32'h00000000;
		12'hcd8:		data <= 32'h00000000;
		12'hcd9:		data <= 32'h00000000;
		12'hcda:		data <= 32'h00000000;
		12'hcdb:		data <= 32'h00000000;
		12'hcdc:		data <= 32'h00000000;
		12'hcdd:		data <= 32'h00000000;
		12'hcde:		data <= 32'h00000000;
		12'hcdf:		data <= 32'h00000000;
		12'hce0:		data <= 32'h00000000;
		12'hce1:		data <= 32'h00000000;
		12'hce2:		data <= 32'h00000000;
		12'hce3:		data <= 32'h00000000;
		12'hce4:		data <= 32'h00000000;
		12'hce5:		data <= 32'h00000000;
		12'hce6:		data <= 32'h00000000;
		12'hce7:		data <= 32'h00000000;
		12'hce8:		data <= 32'h00000000;
		12'hce9:		data <= 32'h00000000;
		12'hcea:		data <= 32'h00000000;
		12'hceb:		data <= 32'h00000000;
		12'hcec:		data <= 32'h00000000;
		12'hced:		data <= 32'h00000000;
		12'hcee:		data <= 32'h00000000;
		12'hcef:		data <= 32'h00000000;
		12'hcf0:		data <= 32'h00000000;
		12'hcf1:		data <= 32'h00000000;
		12'hcf2:		data <= 32'h00000000;
		12'hcf3:		data <= 32'h00000000;
		12'hcf4:		data <= 32'h00000000;
		12'hcf5:		data <= 32'h00000000;
		12'hcf6:		data <= 32'h00000000;
		12'hcf7:		data <= 32'h00000000;
		12'hcf8:		data <= 32'h00000000;
		12'hcf9:		data <= 32'h00000000;
		12'hcfa:		data <= 32'h00000000;
		12'hcfb:		data <= 32'h00000000;
		12'hcfc:		data <= 32'h00000000;
		12'hcfd:		data <= 32'h00000000;
		12'hcfe:		data <= 32'h00000000;
		12'hcff:		data <= 32'h00000000;
		12'hd00:		data <= 32'h00000000;
		12'hd01:		data <= 32'h00000000;
		12'hd02:		data <= 32'h00000000;
		12'hd03:		data <= 32'h00000000;
		12'hd04:		data <= 32'h00000000;
		12'hd05:		data <= 32'h00000000;
		12'hd06:		data <= 32'h00000000;
		12'hd07:		data <= 32'h00000000;
		12'hd08:		data <= 32'h00000000;
		12'hd09:		data <= 32'h00000000;
		12'hd0a:		data <= 32'h00000000;
		12'hd0b:		data <= 32'h00000000;
		12'hd0c:		data <= 32'h00000000;
		12'hd0d:		data <= 32'h00000000;
		12'hd0e:		data <= 32'h00000000;
		12'hd0f:		data <= 32'h00000000;
		12'hd10:		data <= 32'h00000000;
		12'hd11:		data <= 32'h00000000;
		12'hd12:		data <= 32'h00000000;
		12'hd13:		data <= 32'h00000000;
		12'hd14:		data <= 32'h00000000;
		12'hd15:		data <= 32'h00000000;
		12'hd16:		data <= 32'h00000000;
		12'hd17:		data <= 32'h00000000;
		12'hd18:		data <= 32'h00000000;
		12'hd19:		data <= 32'h00000000;
		12'hd1a:		data <= 32'h00000000;
		12'hd1b:		data <= 32'h00000000;
		12'hd1c:		data <= 32'h00000000;
		12'hd1d:		data <= 32'h00000000;
		12'hd1e:		data <= 32'h00000000;
		12'hd1f:		data <= 32'h00000000;
		12'hd20:		data <= 32'h00000000;
		12'hd21:		data <= 32'h00000000;
		12'hd22:		data <= 32'h00000000;
		12'hd23:		data <= 32'h00000000;
		12'hd24:		data <= 32'h00000000;
		12'hd25:		data <= 32'h00000000;
		12'hd26:		data <= 32'h00000000;
		12'hd27:		data <= 32'h00000000;
		12'hd28:		data <= 32'h00000000;
		12'hd29:		data <= 32'h00000000;
		12'hd2a:		data <= 32'h00000000;
		12'hd2b:		data <= 32'h00000000;
		12'hd2c:		data <= 32'h00000000;
		12'hd2d:		data <= 32'h00000000;
		12'hd2e:		data <= 32'h00000000;
		12'hd2f:		data <= 32'h00000000;
		12'hd30:		data <= 32'h00000000;
		12'hd31:		data <= 32'h00000000;
		12'hd32:		data <= 32'h00000000;
		12'hd33:		data <= 32'h00000000;
		12'hd34:		data <= 32'h00000000;
		12'hd35:		data <= 32'h00000000;
		12'hd36:		data <= 32'h00000000;
		12'hd37:		data <= 32'h00000000;
		12'hd38:		data <= 32'h00000000;
		12'hd39:		data <= 32'h00000000;
		12'hd3a:		data <= 32'h00000000;
		12'hd3b:		data <= 32'h00000000;
		12'hd3c:		data <= 32'h00000000;
		12'hd3d:		data <= 32'h00000000;
		12'hd3e:		data <= 32'h00000000;
		12'hd3f:		data <= 32'h00000000;
		12'hd40:		data <= 32'h00000000;
		12'hd41:		data <= 32'h00000000;
		12'hd42:		data <= 32'h00000000;
		12'hd43:		data <= 32'h00000000;
		12'hd44:		data <= 32'h00000000;
		12'hd45:		data <= 32'h00000000;
		12'hd46:		data <= 32'h00000000;
		12'hd47:		data <= 32'h00000000;
		12'hd48:		data <= 32'h00000000;
		12'hd49:		data <= 32'h00000000;
		12'hd4a:		data <= 32'h00000000;
		12'hd4b:		data <= 32'h00000000;
		12'hd4c:		data <= 32'h00000000;
		12'hd4d:		data <= 32'h00000000;
		12'hd4e:		data <= 32'h00000000;
		12'hd4f:		data <= 32'h00000000;
		12'hd50:		data <= 32'h00000000;
		12'hd51:		data <= 32'h00000000;
		12'hd52:		data <= 32'h00000000;
		12'hd53:		data <= 32'h00000000;
		12'hd54:		data <= 32'h00000000;
		12'hd55:		data <= 32'h00000000;
		12'hd56:		data <= 32'h00000000;
		12'hd57:		data <= 32'h00000000;
		12'hd58:		data <= 32'h00000000;
		12'hd59:		data <= 32'h00000000;
		12'hd5a:		data <= 32'h00000000;
		12'hd5b:		data <= 32'h00000000;
		12'hd5c:		data <= 32'h00000000;
		12'hd5d:		data <= 32'h00000000;
		12'hd5e:		data <= 32'h00000000;
		12'hd5f:		data <= 32'h00000000;
		12'hd60:		data <= 32'h00000000;
		12'hd61:		data <= 32'h00000000;
		12'hd62:		data <= 32'h00000000;
		12'hd63:		data <= 32'h00000000;
		12'hd64:		data <= 32'h00000000;
		12'hd65:		data <= 32'h00000000;
		12'hd66:		data <= 32'h00000000;
		12'hd67:		data <= 32'h00000000;
		12'hd68:		data <= 32'h00000000;
		12'hd69:		data <= 32'h00000000;
		12'hd6a:		data <= 32'h00000000;
		12'hd6b:		data <= 32'h00000000;
		12'hd6c:		data <= 32'h00000000;
		12'hd6d:		data <= 32'h00000000;
		12'hd6e:		data <= 32'h00000000;
		12'hd6f:		data <= 32'h00000000;
		12'hd70:		data <= 32'h00000000;
		12'hd71:		data <= 32'h00000000;
		12'hd72:		data <= 32'h00000000;
		12'hd73:		data <= 32'h00000000;
		12'hd74:		data <= 32'h00000000;
		12'hd75:		data <= 32'h00000000;
		12'hd76:		data <= 32'h00000000;
		12'hd77:		data <= 32'h00000000;
		12'hd78:		data <= 32'h00000000;
		12'hd79:		data <= 32'h00000000;
		12'hd7a:		data <= 32'h00000000;
		12'hd7b:		data <= 32'h00000000;
		12'hd7c:		data <= 32'h00000000;
		12'hd7d:		data <= 32'h00000000;
		12'hd7e:		data <= 32'h00000000;
		12'hd7f:		data <= 32'h00000000;
		12'hd80:		data <= 32'h00000000;
		12'hd81:		data <= 32'h00000000;
		12'hd82:		data <= 32'h00000000;
		12'hd83:		data <= 32'h00000000;
		12'hd84:		data <= 32'h00000000;
		12'hd85:		data <= 32'h00000000;
		12'hd86:		data <= 32'h00000000;
		12'hd87:		data <= 32'h00000000;
		12'hd88:		data <= 32'h00000000;
		12'hd89:		data <= 32'h00000000;
		12'hd8a:		data <= 32'h00000000;
		12'hd8b:		data <= 32'h00000000;
		12'hd8c:		data <= 32'h00000000;
		12'hd8d:		data <= 32'h00000000;
		12'hd8e:		data <= 32'h00000000;
		12'hd8f:		data <= 32'h00000000;
		12'hd90:		data <= 32'h00000000;
		12'hd91:		data <= 32'h00000000;
		12'hd92:		data <= 32'h00000000;
		12'hd93:		data <= 32'h00000000;
		12'hd94:		data <= 32'h00000000;
		12'hd95:		data <= 32'h00000000;
		12'hd96:		data <= 32'h00000000;
		12'hd97:		data <= 32'h00000000;
		12'hd98:		data <= 32'h00000000;
		12'hd99:		data <= 32'h00000000;
		12'hd9a:		data <= 32'h00000000;
		12'hd9b:		data <= 32'h00000000;
		12'hd9c:		data <= 32'h00000000;
		12'hd9d:		data <= 32'h00000000;
		12'hd9e:		data <= 32'h00000000;
		12'hd9f:		data <= 32'h00000000;
		12'hda0:		data <= 32'h00000000;
		12'hda1:		data <= 32'h00000000;
		12'hda2:		data <= 32'h00000000;
		12'hda3:		data <= 32'h00000000;
		12'hda4:		data <= 32'h00000000;
		12'hda5:		data <= 32'h00000000;
		12'hda6:		data <= 32'h00000000;
		12'hda7:		data <= 32'h00000000;
		12'hda8:		data <= 32'h00000000;
		12'hda9:		data <= 32'h00000000;
		12'hdaa:		data <= 32'h00000000;
		12'hdab:		data <= 32'h00000000;
		12'hdac:		data <= 32'h00000000;
		12'hdad:		data <= 32'h00000000;
		12'hdae:		data <= 32'h00000000;
		12'hdaf:		data <= 32'h00000000;
		12'hdb0:		data <= 32'h00000000;
		12'hdb1:		data <= 32'h00000000;
		12'hdb2:		data <= 32'h00000000;
		12'hdb3:		data <= 32'h00000000;
		12'hdb4:		data <= 32'h00000000;
		12'hdb5:		data <= 32'h00000000;
		12'hdb6:		data <= 32'h00000000;
		12'hdb7:		data <= 32'h00000000;
		12'hdb8:		data <= 32'h00000000;
		12'hdb9:		data <= 32'h00000000;
		12'hdba:		data <= 32'h00000000;
		12'hdbb:		data <= 32'h00000000;
		12'hdbc:		data <= 32'h00000000;
		12'hdbd:		data <= 32'h00000000;
		12'hdbe:		data <= 32'h00000000;
		12'hdbf:		data <= 32'h00000000;
		12'hdc0:		data <= 32'h00000000;
		12'hdc1:		data <= 32'h00000000;
		12'hdc2:		data <= 32'h00000000;
		12'hdc3:		data <= 32'h00000000;
		12'hdc4:		data <= 32'h00000000;
		12'hdc5:		data <= 32'h00000000;
		12'hdc6:		data <= 32'h00000000;
		12'hdc7:		data <= 32'h00000000;
		12'hdc8:		data <= 32'h00000000;
		12'hdc9:		data <= 32'h00000000;
		12'hdca:		data <= 32'h00000000;
		12'hdcb:		data <= 32'h00000000;
		12'hdcc:		data <= 32'h00000000;
		12'hdcd:		data <= 32'h00000000;
		12'hdce:		data <= 32'h00000000;
		12'hdcf:		data <= 32'h00000000;
		12'hdd0:		data <= 32'h00000000;
		12'hdd1:		data <= 32'h00000000;
		12'hdd2:		data <= 32'h00000000;
		12'hdd3:		data <= 32'h00000000;
		12'hdd4:		data <= 32'h00000000;
		12'hdd5:		data <= 32'h00000000;
		12'hdd6:		data <= 32'h00000000;
		12'hdd7:		data <= 32'h00000000;
		12'hdd8:		data <= 32'h00000000;
		12'hdd9:		data <= 32'h00000000;
		12'hdda:		data <= 32'h00000000;
		12'hddb:		data <= 32'h00000000;
		12'hddc:		data <= 32'h00000000;
		12'hddd:		data <= 32'h00000000;
		12'hdde:		data <= 32'h00000000;
		12'hddf:		data <= 32'h00000000;
		12'hde0:		data <= 32'h00000000;
		12'hde1:		data <= 32'h00000000;
		12'hde2:		data <= 32'h00000000;
		12'hde3:		data <= 32'h00000000;
		12'hde4:		data <= 32'h00000000;
		12'hde5:		data <= 32'h00000000;
		12'hde6:		data <= 32'h00000000;
		12'hde7:		data <= 32'h00000000;
		12'hde8:		data <= 32'h00000000;
		12'hde9:		data <= 32'h00000000;
		12'hdea:		data <= 32'h00000000;
		12'hdeb:		data <= 32'h00000000;
		12'hdec:		data <= 32'h00000000;
		12'hded:		data <= 32'h00000000;
		12'hdee:		data <= 32'h00000000;
		12'hdef:		data <= 32'h00000000;
		12'hdf0:		data <= 32'h00000000;
		12'hdf1:		data <= 32'h00000000;
		12'hdf2:		data <= 32'h00000000;
		12'hdf3:		data <= 32'h00000000;
		12'hdf4:		data <= 32'h00000000;
		12'hdf5:		data <= 32'h00000000;
		12'hdf6:		data <= 32'h00000000;
		12'hdf7:		data <= 32'h00000000;
		12'hdf8:		data <= 32'h00000000;
		12'hdf9:		data <= 32'h00000000;
		12'hdfa:		data <= 32'h00000000;
		12'hdfb:		data <= 32'h00000000;
		12'hdfc:		data <= 32'h00000000;
		12'hdfd:		data <= 32'h00000000;
		12'hdfe:		data <= 32'h00000000;
		12'hdff:		data <= 32'h00000000;
		12'he00:		data <= 32'h00000000;
		12'he01:		data <= 32'h00000000;
		12'he02:		data <= 32'h00000000;
		12'he03:		data <= 32'h00000000;
		12'he04:		data <= 32'h00000000;
		12'he05:		data <= 32'h00000000;
		12'he06:		data <= 32'h00000000;
		12'he07:		data <= 32'h00000000;
		12'he08:		data <= 32'h00000000;
		12'he09:		data <= 32'h00000000;
		12'he0a:		data <= 32'h00000000;
		12'he0b:		data <= 32'h00000000;
		12'he0c:		data <= 32'h00000000;
		12'he0d:		data <= 32'h00000000;
		12'he0e:		data <= 32'h00000000;
		12'he0f:		data <= 32'h00000000;
		12'he10:		data <= 32'h00000000;
		12'he11:		data <= 32'h00000000;
		12'he12:		data <= 32'h00000000;
		12'he13:		data <= 32'h00000000;
		12'he14:		data <= 32'h00000000;
		12'he15:		data <= 32'h00000000;
		12'he16:		data <= 32'h00000000;
		12'he17:		data <= 32'h00000000;
		12'he18:		data <= 32'h00000000;
		12'he19:		data <= 32'h00000000;
		12'he1a:		data <= 32'h00000000;
		12'he1b:		data <= 32'h00000000;
		12'he1c:		data <= 32'h00000000;
		12'he1d:		data <= 32'h00000000;
		12'he1e:		data <= 32'h00000000;
		12'he1f:		data <= 32'h00000000;
		12'he20:		data <= 32'h00000000;
		12'he21:		data <= 32'h00000000;
		12'he22:		data <= 32'h00000000;
		12'he23:		data <= 32'h00000000;
		12'he24:		data <= 32'h00000000;
		12'he25:		data <= 32'h00000000;
		12'he26:		data <= 32'h00000000;
		12'he27:		data <= 32'h00000000;
		12'he28:		data <= 32'h00000000;
		12'he29:		data <= 32'h00000000;
		12'he2a:		data <= 32'h00000000;
		12'he2b:		data <= 32'h00000000;
		12'he2c:		data <= 32'h00000000;
		12'he2d:		data <= 32'h00000000;
		12'he2e:		data <= 32'h00000000;
		12'he2f:		data <= 32'h00000000;
		12'he30:		data <= 32'h00000000;
		12'he31:		data <= 32'h00000000;
		12'he32:		data <= 32'h00000000;
		12'he33:		data <= 32'h00000000;
		12'he34:		data <= 32'h00000000;
		12'he35:		data <= 32'h00000000;
		12'he36:		data <= 32'h00000000;
		12'he37:		data <= 32'h00000000;
		12'he38:		data <= 32'h00000000;
		12'he39:		data <= 32'h00000000;
		12'he3a:		data <= 32'h00000000;
		12'he3b:		data <= 32'h00000000;
		12'he3c:		data <= 32'h00000000;
		12'he3d:		data <= 32'h00000000;
		12'he3e:		data <= 32'h00000000;
		12'he3f:		data <= 32'h00000000;
		12'he40:		data <= 32'h00000000;
		12'he41:		data <= 32'h00000000;
		12'he42:		data <= 32'h00000000;
		12'he43:		data <= 32'h00000000;
		12'he44:		data <= 32'h00000000;
		12'he45:		data <= 32'h00000000;
		12'he46:		data <= 32'h00000000;
		12'he47:		data <= 32'h00000000;
		12'he48:		data <= 32'h00000000;
		12'he49:		data <= 32'h00000000;
		12'he4a:		data <= 32'h00000000;
		12'he4b:		data <= 32'h00000000;
		12'he4c:		data <= 32'h00000000;
		12'he4d:		data <= 32'h00000000;
		12'he4e:		data <= 32'h00000000;
		12'he4f:		data <= 32'h00000000;
		12'he50:		data <= 32'h00000000;
		12'he51:		data <= 32'h00000000;
		12'he52:		data <= 32'h00000000;
		12'he53:		data <= 32'h00000000;
		12'he54:		data <= 32'h00000000;
		12'he55:		data <= 32'h00000000;
		12'he56:		data <= 32'h00000000;
		12'he57:		data <= 32'h00000000;
		12'he58:		data <= 32'h00000000;
		12'he59:		data <= 32'h00000000;
		12'he5a:		data <= 32'h00000000;
		12'he5b:		data <= 32'h00000000;
		12'he5c:		data <= 32'h00000000;
		12'he5d:		data <= 32'h00000000;
		12'he5e:		data <= 32'h00000000;
		12'he5f:		data <= 32'h00000000;
		12'he60:		data <= 32'h00000000;
		12'he61:		data <= 32'h00000000;
		12'he62:		data <= 32'h00000000;
		12'he63:		data <= 32'h00000000;
		12'he64:		data <= 32'h00000000;
		12'he65:		data <= 32'h00000000;
		12'he66:		data <= 32'h00000000;
		12'he67:		data <= 32'h00000000;
		12'he68:		data <= 32'h00000000;
		12'he69:		data <= 32'h00000000;
		12'he6a:		data <= 32'h00000000;
		12'he6b:		data <= 32'h00000000;
		12'he6c:		data <= 32'h00000000;
		12'he6d:		data <= 32'h00000000;
		12'he6e:		data <= 32'h00000000;
		12'he6f:		data <= 32'h00000000;
		12'he70:		data <= 32'h00000000;
		12'he71:		data <= 32'h00000000;
		12'he72:		data <= 32'h00000000;
		12'he73:		data <= 32'h00000000;
		12'he74:		data <= 32'h00000000;
		12'he75:		data <= 32'h00000000;
		12'he76:		data <= 32'h00000000;
		12'he77:		data <= 32'h00000000;
		12'he78:		data <= 32'h00000000;
		12'he79:		data <= 32'h00000000;
		12'he7a:		data <= 32'h00000000;
		12'he7b:		data <= 32'h00000000;
		12'he7c:		data <= 32'h00000000;
		12'he7d:		data <= 32'h00000000;
		12'he7e:		data <= 32'h00000000;
		12'he7f:		data <= 32'h00000000;
		12'he80:		data <= 32'h00000000;
		12'he81:		data <= 32'h00000000;
		12'he82:		data <= 32'h00000000;
		12'he83:		data <= 32'h00000000;
		12'he84:		data <= 32'h00000000;
		12'he85:		data <= 32'h00000000;
		12'he86:		data <= 32'h00000000;
		12'he87:		data <= 32'h00000000;
		12'he88:		data <= 32'h00000000;
		12'he89:		data <= 32'h00000000;
		12'he8a:		data <= 32'h00000000;
		12'he8b:		data <= 32'h00000000;
		12'he8c:		data <= 32'h00000000;
		12'he8d:		data <= 32'h00000000;
		12'he8e:		data <= 32'h00000000;
		12'he8f:		data <= 32'h00000000;
		12'he90:		data <= 32'h00000000;
		12'he91:		data <= 32'h00000000;
		12'he92:		data <= 32'h00000000;
		12'he93:		data <= 32'h00000000;
		12'he94:		data <= 32'h00000000;
		12'he95:		data <= 32'h00000000;
		12'he96:		data <= 32'h00000000;
		12'he97:		data <= 32'h00000000;
		12'he98:		data <= 32'h00000000;
		12'he99:		data <= 32'h00000000;
		12'he9a:		data <= 32'h00000000;
		12'he9b:		data <= 32'h00000000;
		12'he9c:		data <= 32'h00000000;
		12'he9d:		data <= 32'h00000000;
		12'he9e:		data <= 32'h00000000;
		12'he9f:		data <= 32'h00000000;
		12'hea0:		data <= 32'h00000000;
		12'hea1:		data <= 32'h00000000;
		12'hea2:		data <= 32'h00000000;
		12'hea3:		data <= 32'h00000000;
		12'hea4:		data <= 32'h00000000;
		12'hea5:		data <= 32'h00000000;
		12'hea6:		data <= 32'h00000000;
		12'hea7:		data <= 32'h00000000;
		12'hea8:		data <= 32'h00000000;
		12'hea9:		data <= 32'h00000000;
		12'heaa:		data <= 32'h00000000;
		12'heab:		data <= 32'h00000000;
		12'heac:		data <= 32'h00000000;
		12'head:		data <= 32'h00000000;
		12'heae:		data <= 32'h00000000;
		12'heaf:		data <= 32'h00000000;
		12'heb0:		data <= 32'h00000000;
		12'heb1:		data <= 32'h00000000;
		12'heb2:		data <= 32'h00000000;
		12'heb3:		data <= 32'h00000000;
		12'heb4:		data <= 32'h00000000;
		12'heb5:		data <= 32'h00000000;
		12'heb6:		data <= 32'h00000000;
		12'heb7:		data <= 32'h00000000;
		12'heb8:		data <= 32'h00000000;
		12'heb9:		data <= 32'h00000000;
		12'heba:		data <= 32'h00000000;
		12'hebb:		data <= 32'h00000000;
		12'hebc:		data <= 32'h00000000;
		12'hebd:		data <= 32'h00000000;
		12'hebe:		data <= 32'h00000000;
		12'hebf:		data <= 32'h00000000;
		12'hec0:		data <= 32'h00000000;
		12'hec1:		data <= 32'h00000000;
		12'hec2:		data <= 32'h00000000;
		12'hec3:		data <= 32'h00000000;
		12'hec4:		data <= 32'h00000000;
		12'hec5:		data <= 32'h00000000;
		12'hec6:		data <= 32'h00000000;
		12'hec7:		data <= 32'h00000000;
		12'hec8:		data <= 32'h00000000;
		12'hec9:		data <= 32'h00000000;
		12'heca:		data <= 32'h00000000;
		12'hecb:		data <= 32'h00000000;
		12'hecc:		data <= 32'h00000000;
		12'hecd:		data <= 32'h00000000;
		12'hece:		data <= 32'h00000000;
		12'hecf:		data <= 32'h00000000;
		12'hed0:		data <= 32'h00000000;
		12'hed1:		data <= 32'h00000000;
		12'hed2:		data <= 32'h00000000;
		12'hed3:		data <= 32'h00000000;
		12'hed4:		data <= 32'h00000000;
		12'hed5:		data <= 32'h00000000;
		12'hed6:		data <= 32'h00000000;
		12'hed7:		data <= 32'h00000000;
		12'hed8:		data <= 32'h00000000;
		12'hed9:		data <= 32'h00000000;
		12'heda:		data <= 32'h00000000;
		12'hedb:		data <= 32'h00000000;
		12'hedc:		data <= 32'h00000000;
		12'hedd:		data <= 32'h00000000;
		12'hede:		data <= 32'h00000000;
		12'hedf:		data <= 32'h00000000;
		12'hee0:		data <= 32'h00000000;
		12'hee1:		data <= 32'h00000000;
		12'hee2:		data <= 32'h00000000;
		12'hee3:		data <= 32'h00000000;
		12'hee4:		data <= 32'h00000000;
		12'hee5:		data <= 32'h00000000;
		12'hee6:		data <= 32'h00000000;
		12'hee7:		data <= 32'h00000000;
		12'hee8:		data <= 32'h00000000;
		12'hee9:		data <= 32'h00000000;
		12'heea:		data <= 32'h00000000;
		12'heeb:		data <= 32'h00000000;
		12'heec:		data <= 32'h00000000;
		12'heed:		data <= 32'h00000000;
		12'heee:		data <= 32'h00000000;
		12'heef:		data <= 32'h00000000;
		12'hef0:		data <= 32'h00000000;
		12'hef1:		data <= 32'h00000000;
		12'hef2:		data <= 32'h00000000;
		12'hef3:		data <= 32'h00000000;
		12'hef4:		data <= 32'h00000000;
		12'hef5:		data <= 32'h00000000;
		12'hef6:		data <= 32'h00000000;
		12'hef7:		data <= 32'h00000000;
		12'hef8:		data <= 32'h00000000;
		12'hef9:		data <= 32'h00000000;
		12'hefa:		data <= 32'h00000000;
		12'hefb:		data <= 32'h00000000;
		12'hefc:		data <= 32'h00000000;
		12'hefd:		data <= 32'h00000000;
		12'hefe:		data <= 32'h00000000;
		12'heff:		data <= 32'h00000000;
		12'hf00:		data <= 32'h00000000;
		12'hf01:		data <= 32'h00000000;
		12'hf02:		data <= 32'h00000000;
		12'hf03:		data <= 32'h00000000;
		12'hf04:		data <= 32'h00000000;
		12'hf05:		data <= 32'h00000000;
		12'hf06:		data <= 32'h00000000;
		12'hf07:		data <= 32'h00000000;
		12'hf08:		data <= 32'h00000000;
		12'hf09:		data <= 32'h00000000;
		12'hf0a:		data <= 32'h00000000;
		12'hf0b:		data <= 32'h00000000;
		12'hf0c:		data <= 32'h00000000;
		12'hf0d:		data <= 32'h00000000;
		12'hf0e:		data <= 32'h00000000;
		12'hf0f:		data <= 32'h00000000;
		12'hf10:		data <= 32'h00000000;
		12'hf11:		data <= 32'h00000000;
		12'hf12:		data <= 32'h00000000;
		12'hf13:		data <= 32'h00000000;
		12'hf14:		data <= 32'h00000000;
		12'hf15:		data <= 32'h00000000;
		12'hf16:		data <= 32'h00000000;
		12'hf17:		data <= 32'h00000000;
		12'hf18:		data <= 32'h00000000;
		12'hf19:		data <= 32'h00000000;
		12'hf1a:		data <= 32'h00000000;
		12'hf1b:		data <= 32'h00000000;
		12'hf1c:		data <= 32'h00000000;
		12'hf1d:		data <= 32'h00000000;
		12'hf1e:		data <= 32'h00000000;
		12'hf1f:		data <= 32'h00000000;
		12'hf20:		data <= 32'h00000000;
		12'hf21:		data <= 32'h00000000;
		12'hf22:		data <= 32'h00000000;
		12'hf23:		data <= 32'h00000000;
		12'hf24:		data <= 32'h00000000;
		12'hf25:		data <= 32'h00000000;
		12'hf26:		data <= 32'h00000000;
		12'hf27:		data <= 32'h00000000;
		12'hf28:		data <= 32'h00000000;
		12'hf29:		data <= 32'h00000000;
		12'hf2a:		data <= 32'h00000000;
		12'hf2b:		data <= 32'h00000000;
		12'hf2c:		data <= 32'h00000000;
		12'hf2d:		data <= 32'h00000000;
		12'hf2e:		data <= 32'h00000000;
		12'hf2f:		data <= 32'h00000000;
		12'hf30:		data <= 32'h00000000;
		12'hf31:		data <= 32'h00000000;
		12'hf32:		data <= 32'h00000000;
		12'hf33:		data <= 32'h00000000;
		12'hf34:		data <= 32'h00000000;
		12'hf35:		data <= 32'h00000000;
		12'hf36:		data <= 32'h00000000;
		12'hf37:		data <= 32'h00000000;
		12'hf38:		data <= 32'h00000000;
		12'hf39:		data <= 32'h00000000;
		12'hf3a:		data <= 32'h00000000;
		12'hf3b:		data <= 32'h00000000;
		12'hf3c:		data <= 32'h00000000;
		12'hf3d:		data <= 32'h00000000;
		12'hf3e:		data <= 32'h00000000;
		12'hf3f:		data <= 32'h00000000;
		12'hf40:		data <= 32'h00000000;
		12'hf41:		data <= 32'h00000000;
		12'hf42:		data <= 32'h00000000;
		12'hf43:		data <= 32'h00000000;
		12'hf44:		data <= 32'h00000000;
		12'hf45:		data <= 32'h00000000;
		12'hf46:		data <= 32'h00000000;
		12'hf47:		data <= 32'h00000000;
		12'hf48:		data <= 32'h00000000;
		12'hf49:		data <= 32'h00000000;
		12'hf4a:		data <= 32'h00000000;
		12'hf4b:		data <= 32'h00000000;
		12'hf4c:		data <= 32'h00000000;
		12'hf4d:		data <= 32'h00000000;
		12'hf4e:		data <= 32'h00000000;
		12'hf4f:		data <= 32'h00000000;
		12'hf50:		data <= 32'h00000000;
		12'hf51:		data <= 32'h00000000;
		12'hf52:		data <= 32'h00000000;
		12'hf53:		data <= 32'h00000000;
		12'hf54:		data <= 32'h00000000;
		12'hf55:		data <= 32'h00000000;
		12'hf56:		data <= 32'h00000000;
		12'hf57:		data <= 32'h00000000;
		12'hf58:		data <= 32'h00000000;
		12'hf59:		data <= 32'h00000000;
		12'hf5a:		data <= 32'h00000000;
		12'hf5b:		data <= 32'h00000000;
		12'hf5c:		data <= 32'h00000000;
		12'hf5d:		data <= 32'h00000000;
		12'hf5e:		data <= 32'h00000000;
		12'hf5f:		data <= 32'h00000000;
		12'hf60:		data <= 32'h00000000;
		12'hf61:		data <= 32'h00000000;
		12'hf62:		data <= 32'h00000000;
		12'hf63:		data <= 32'h00000000;
		12'hf64:		data <= 32'h00000000;
		12'hf65:		data <= 32'h00000000;
		12'hf66:		data <= 32'h00000000;
		12'hf67:		data <= 32'h00000000;
		12'hf68:		data <= 32'h00000000;
		12'hf69:		data <= 32'h00000000;
		12'hf6a:		data <= 32'h00000000;
		12'hf6b:		data <= 32'h00000000;
		12'hf6c:		data <= 32'h00000000;
		12'hf6d:		data <= 32'h00000000;
		12'hf6e:		data <= 32'h00000000;
		12'hf6f:		data <= 32'h00000000;
		12'hf70:		data <= 32'h00000000;
		12'hf71:		data <= 32'h00000000;
		12'hf72:		data <= 32'h00000000;
		12'hf73:		data <= 32'h00000000;
		12'hf74:		data <= 32'h00000000;
		12'hf75:		data <= 32'h00000000;
		12'hf76:		data <= 32'h00000000;
		12'hf77:		data <= 32'h00000000;
		12'hf78:		data <= 32'h00000000;
		12'hf79:		data <= 32'h00000000;
		12'hf7a:		data <= 32'h00000000;
		12'hf7b:		data <= 32'h00000000;
		12'hf7c:		data <= 32'h00000000;
		12'hf7d:		data <= 32'h00000000;
		12'hf7e:		data <= 32'h00000000;
		12'hf7f:		data <= 32'h00000000;
		12'hf80:		data <= 32'h00000000;
		12'hf81:		data <= 32'h00000000;
		12'hf82:		data <= 32'h00000000;
		12'hf83:		data <= 32'h00000000;
		12'hf84:		data <= 32'h00000000;
		12'hf85:		data <= 32'h00000000;
		12'hf86:		data <= 32'h00000000;
		12'hf87:		data <= 32'h00000000;
		12'hf88:		data <= 32'h00000000;
		12'hf89:		data <= 32'h00000000;
		12'hf8a:		data <= 32'h00000000;
		12'hf8b:		data <= 32'h00000000;
		12'hf8c:		data <= 32'h00000000;
		12'hf8d:		data <= 32'h00000000;
		12'hf8e:		data <= 32'h00000000;
		12'hf8f:		data <= 32'h00000000;
		12'hf90:		data <= 32'h00000000;
		12'hf91:		data <= 32'h00000000;
		12'hf92:		data <= 32'h00000000;
		12'hf93:		data <= 32'h00000000;
		12'hf94:		data <= 32'h00000000;
		12'hf95:		data <= 32'h00000000;
		12'hf96:		data <= 32'h00000000;
		12'hf97:		data <= 32'h00000000;
		12'hf98:		data <= 32'h00000000;
		12'hf99:		data <= 32'h00000000;
		12'hf9a:		data <= 32'h00000000;
		12'hf9b:		data <= 32'h00000000;
		12'hf9c:		data <= 32'h00000000;
		12'hf9d:		data <= 32'h00000000;
		12'hf9e:		data <= 32'h00000000;
		12'hf9f:		data <= 32'h00000000;
		12'hfa0:		data <= 32'h00000000;
		12'hfa1:		data <= 32'h00000000;
		12'hfa2:		data <= 32'h00000000;
		12'hfa3:		data <= 32'h00000000;
		12'hfa4:		data <= 32'h00000000;
		12'hfa5:		data <= 32'h00000000;
		12'hfa6:		data <= 32'h00000000;
		12'hfa7:		data <= 32'h00000000;
		12'hfa8:		data <= 32'h00000000;
		12'hfa9:		data <= 32'h00000000;
		12'hfaa:		data <= 32'h00000000;
		12'hfab:		data <= 32'h00000000;
		12'hfac:		data <= 32'h00000000;
		12'hfad:		data <= 32'h00000000;
		12'hfae:		data <= 32'h00000000;
		12'hfaf:		data <= 32'h00000000;
		12'hfb0:		data <= 32'h00000000;
		12'hfb1:		data <= 32'h00000000;
		12'hfb2:		data <= 32'h00000000;
		12'hfb3:		data <= 32'h00000000;
		12'hfb4:		data <= 32'h00000000;
		12'hfb5:		data <= 32'h00000000;
		12'hfb6:		data <= 32'h00000000;
		12'hfb7:		data <= 32'h00000000;
		12'hfb8:		data <= 32'h00000000;
		12'hfb9:		data <= 32'h00000000;
		12'hfba:		data <= 32'h00000000;
		12'hfbb:		data <= 32'h00000000;
		12'hfbc:		data <= 32'h00000000;
		12'hfbd:		data <= 32'h00000000;
		12'hfbe:		data <= 32'h00000000;
		12'hfbf:		data <= 32'h00000000;
		12'hfc0:		data <= 32'h00000000;
		12'hfc1:		data <= 32'h00000000;
		12'hfc2:		data <= 32'h00000000;
		12'hfc3:		data <= 32'h00000000;
		12'hfc4:		data <= 32'h00000000;
		12'hfc5:		data <= 32'h00000000;
		12'hfc6:		data <= 32'h00000000;
		12'hfc7:		data <= 32'h00000000;
		12'hfc8:		data <= 32'h00000000;
		12'hfc9:		data <= 32'h00000000;
		12'hfca:		data <= 32'h00000000;
		12'hfcb:		data <= 32'h00000000;
		12'hfcc:		data <= 32'h00000000;
		12'hfcd:		data <= 32'h00000000;
		12'hfce:		data <= 32'h00000000;
		12'hfcf:		data <= 32'h00000000;
		12'hfd0:		data <= 32'h00000000;
		12'hfd1:		data <= 32'h00000000;
		12'hfd2:		data <= 32'h00000000;
		12'hfd3:		data <= 32'h00000000;
		12'hfd4:		data <= 32'h00000000;
		12'hfd5:		data <= 32'h00000000;
		12'hfd6:		data <= 32'h00000000;
		12'hfd7:		data <= 32'h00000000;
		12'hfd8:		data <= 32'h00000000;
		12'hfd9:		data <= 32'h00000000;
		12'hfda:		data <= 32'h00000000;
		12'hfdb:		data <= 32'h00000000;
		12'hfdc:		data <= 32'h00000000;
		12'hfdd:		data <= 32'h00000000;
		12'hfde:		data <= 32'h00000000;
		12'hfdf:		data <= 32'h00000000;
		12'hfe0:		data <= 32'h00000000;
		12'hfe1:		data <= 32'h00000000;
		12'hfe2:		data <= 32'h00000000;
		12'hfe3:		data <= 32'h00000000;
		12'hfe4:		data <= 32'h00000000;
		12'hfe5:		data <= 32'h00000000;
		12'hfe6:		data <= 32'h00000000;
		12'hfe7:		data <= 32'h00000000;
		12'hfe8:		data <= 32'h00000000;
		12'hfe9:		data <= 32'h00000000;
		12'hfea:		data <= 32'h00000000;
		12'hfeb:		data <= 32'h00000000;
		12'hfec:		data <= 32'h00000000;
		12'hfed:		data <= 32'h00000000;
		12'hfee:		data <= 32'h00000000;
		12'hfef:		data <= 32'h00000000;
		12'hff0:		data <= 32'h00000000;
		12'hff1:		data <= 32'h00000000;
		12'hff2:		data <= 32'h00000000;
		12'hff3:		data <= 32'h00000000;
		12'hff4:		data <= 32'h00000000;
		12'hff5:		data <= 32'h00000000;
		12'hff6:		data <= 32'h00000000;
		12'hff7:		data <= 32'h00000000;
		12'hff8:		data <= 32'h00000000;
		12'hff9:		data <= 32'h00000000;
		12'hffa:		data <= 32'h00000000;
		12'hffb:		data <= 32'h00000000;
		12'hffc:		data <= 32'h00000000;
		12'hffd:		data <= 32'h00000000;
		12'hffe:		data <= 32'h00000000;
		12'hfff:		data <= 32'h00000000;
		default:	data <= 32'hf0000000;
		endcase
	end
	
endmodule
