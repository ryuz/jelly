
`default_nettype none

module clkgen_clkdiv
        (
            input   var logic   reset_n,
            input   var logic   clk_in,
            output  var logic   clk_out
        );

endmodule


`default_nettype wire


