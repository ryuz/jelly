module Gowin_PLL_dvi_vga(
    clkin,
    init_clk,
    clkout0,
    clkout1,
    lock
);

input clkin;
input init_clk;
output clkout0;
output clkout1;
output lock;

endmodule
