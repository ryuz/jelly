
`timescale 1ns / 1ps
`default_nettype none


module OSER10
        (
            output  var logic   Q     ,
            input   var logic   D0    ,
            input   var logic   D1    ,
            input   var logic   D2    ,
            input   var logic   D3    ,
            input   var logic   D4    ,
            input   var logic   D5    ,
            input   var logic   D6    ,
            input   var logic   D7    ,
            input   var logic   D8    ,
            input   var logic   D9    ,
            input   var logic   PCLK  ,
            input   var logic   FCLK  ,
            input   var logic   RESET 
        );
    
endmodule


`default_nettype wire


