
`timescale 1ns / 1ps
`default_nettype none


module tb_top();
    
    initial begin
        $dumpfile("tb_top.vcd");
        $dumpvars(0, tb_top);
    
    #40000000
        $finish;
    end
    

    // -----------------------------
    //  reset & clock
    // -----------------------------

    localparam RATE100 = 1000.0/100.00;
    localparam RATE200 = 1000.0/200.00;
    localparam RATE250 = 1000.0/250.00;
    localparam RATE133 = 1000.0/133.33;

    reg			reset = 1;
    initial #100 reset = 0;

    reg			clk100 = 1'b1;
    always #(RATE100/2.0) clk100 <= ~clk100;

    reg			clk200 = 1'b1;
    always #(RATE200/2.0) clk200 <= ~clk200;

    reg			clk250 = 1'b1;
    always #(RATE250/2.0) clk250 <= ~clk250;


    // -----------------------------
    //  target
    // -----------------------------

    parameter   int     WIDTH_BITS  = 16;
    parameter   int     HEIGHT_BITS = 16;
    parameter   int     IMG_WIDTH   = 3280 / 2;
    parameter   int     IMG_HEIGHT  = 2464 / 2;

    kv260_imx219
            #(
                .WIDTH_BITS     (WIDTH_BITS     ),
                .HEIGHT_BITS    (HEIGHT_BITS    ),
                .IMG_WIDTH      (IMG_WIDTH      ),
                .IMG_HEIGHT     (IMG_HEIGHT     )
            )
        i_top
            (
                .cam_clk_p      (),
                .cam_clk_n      (),
                .cam_data_p     (),
                .cam_data_n     (),
                .cam_scl        (),
                .cam_sda        (),
                .cam_enable     (),
                .fan_en         (),
                .pmod           ()
            );
    

    // -----------------------------
    //  Clock & Reset
    // -----------------------------
    
    always_comb force i_top.i_design_1.reset  = reset;
    always_comb force i_top.i_design_1.clk100 = clk100;
    always_comb force i_top.i_design_1.clk200 = clk200;
    always_comb force i_top.i_design_1.clk250 = clk250;

    always_comb force i_top.i_design_1.m_axi4l_peri_aresetn = ~reset;
    always_comb force i_top.i_design_1.m_axi4l_peri_aclk    = clk250;

    always_comb force i_top.i_design_1.s_axi4_mem_aresetn = ~reset;
    always_comb force i_top.i_design_1.s_axi4_mem_aclk    = clk250;
    

    // -----------------------------
    //  Video input
    // -----------------------------

    logic   axi4s_src_aresetn;
    logic   axi4s_src_aclk;

    assign axi4s_src_aresetn = i_top.i_mipi_csi2_rx.m_axi4s_aresetn;
    assign axi4s_src_aclk    = i_top.i_mipi_csi2_rx.m_axi4s_aclk;

    jelly3_axi4s_if
            #(
                .USER_BITS      (1),
                .DATA_BITS      (10)
            )
        i_axi4s_src
            (
                .aresetn        (axi4s_src_aresetn),
                .aclk           (axi4s_src_aclk)
            );
    
    always_comb force i_top.i_mipi_csi2_rx.axi4s_tuser  = i_axi4s_src.tuser ;
    always_comb force i_top.i_mipi_csi2_rx.axi4s_tlast  = i_axi4s_src.tlast ;
    always_comb force i_top.i_mipi_csi2_rx.axi4s_tdata  = i_axi4s_src.tdata ;
    always_comb force i_top.i_mipi_csi2_rx.axi4s_tvalid = i_axi4s_src.tvalid;
    assign i_axi4s_src.tready = i_top.i_mipi_csi2_rx.axi4s_tready;


    localparam  SIM_IMG_WIDTH  = 256;
    localparam  SIM_IMG_HEIGHT = 256;

    // master
    jelly3_model_axi4s_m
            #(
                .IMG_WIDTH          (SIM_IMG_WIDTH),
                .IMG_HEIGHT         (SIM_IMG_HEIGHT),
                .FILE_NAME          (),//"../Mandrill_256x256.ppm"),
                .FILE_IMG_WIDTH     (256),
                .FILE_IMG_HEIGHT    (256),
                .BUSY_RATE          (0),
                .RANDOM_SEED        (0)
            )
        u_model_axi4s_m
            (
                .aclken             (1'b1           ),
                .enable             (1'b1           ),
                .busy               (               ),

                .m_axi4s            (i_axi4s_src.m  ),
                .out_x              (               ),
                .out_y              (               ),
                .out_f              (               )
            );


    // -----------------------------
    //  Peripheral Bus
    // -----------------------------

    logic   [0:0]   axi4l_peri_aresetn  ;
    logic           axi4l_peri_aclk     ;

    jelly3_axi4l_if
            #(
                .ADDR_BITS  (40                     ),
                .DATA_BITS  (64                     )
            )
        axi4l_peri
            (
                .aresetn    (axi4l_peri_aresetn     ),
                .aclk       (axi4l_peri_aclk        )
            );

    /*
    logic   [39:0]  axi4l_peri_araddr   ;
    logic   [2:0]   axi4l_peri_arprot   ;
    logic           axi4l_peri_arready  ;
    logic           axi4l_peri_arvalid  ;
    logic   [39:0]  axi4l_peri_awaddr   ;
    logic   [2:0]   axi4l_peri_awprot   ;
    logic           axi4l_peri_awready  ;
    logic           axi4l_peri_awvalid  ;
    logic           axi4l_peri_bready   ;
    logic   [1:0]   axi4l_peri_bresp    ;
    logic           axi4l_peri_bvalid   ;
    logic   [63:0]  axi4l_peri_rdata    ;
    logic           axi4l_peri_rready   ;
    logic   [1:0]   axi4l_peri_rresp    ;
    logic           axi4l_peri_rvalid   ;
    logic   [63:0]  axi4l_peri_wdata    ;
    logic           axi4l_peri_wready   ;
    logic   [7:0]   axi4l_peri_wstrb    ;
    logic           axi4l_peri_wvalid   ;
    */

    assign axi4l_peri_aresetn = i_top.i_design_1.axi4l_peri_aresetn ;
    assign axi4l_peri_aclk    = i_top.i_design_1.axi4l_peri_aclk    ;

    assign axi4l_peri.awready = i_top.i_design_1.axi4l_peri_awready ;
    assign axi4l_peri.wready  = i_top.i_design_1.axi4l_peri_wready  ;
    assign axi4l_peri.bready  = i_top.i_design_1.axi4l_peri_bready  ;
    assign axi4l_peri.bresp   = i_top.i_design_1.axi4l_peri_bresp   ;
    assign axi4l_peri.bvalid  = i_top.i_design_1.axi4l_peri_bvalid  ;
    assign axi4l_peri.arready = i_top.i_design_1.axi4l_peri_arready ;
    assign axi4l_peri.rdata   = i_top.i_design_1.axi4l_peri_rdata   ;
    assign axi4l_peri.rresp   = i_top.i_design_1.axi4l_peri_rresp   ;
    assign axi4l_peri.rvalid  = i_top.i_design_1.axi4l_peri_rvalid  ;

    always_comb force i_top.i_design_1.axi4l_peri_awaddr  = axi4l_peri.awaddr ;
    always_comb force i_top.i_design_1.axi4l_peri_awprot  = axi4l_peri.awprot ;
    always_comb force i_top.i_design_1.axi4l_peri_awvalid = axi4l_peri.awvalid;
    always_comb force i_top.i_design_1.axi4l_peri_wdata   = axi4l_peri.wdata  ;
    always_comb force i_top.i_design_1.axi4l_peri_wstrb   = axi4l_peri.wstrb  ;
    always_comb force i_top.i_design_1.axi4l_peri_wvalid  = axi4l_peri.wvalid ;
    always_comb force i_top.i_design_1.axi4l_peri_bready  = axi4l_peri.bready ;
    always_comb force i_top.i_design_1.axi4l_peri_araddr  = axi4l_peri.araddr ;
    always_comb force i_top.i_design_1.axi4l_peri_arprot  = axi4l_peri.arprot ;
    always_comb force i_top.i_design_1.axi4l_peri_arvalid = axi4l_peri.arvalid;
    always_comb force i_top.i_design_1.axi4l_peri_rready  = axi4l_peri.rready ;




    // -----------------------------
    //  access
    // -----------------------------

    
    localparam type axi4l_addr_t = logic [axi4l_peri.ADDR_BITS-1:0];
    localparam type axi4l_data_t = logic [axi4l_peri.DATA_BITS-1:0];

    localparam  axi4l_addr_t    ADR_GPIO = axi4l_addr_t'(40'ha000_0000);
    localparam  axi4l_addr_t    ADR_FMTR = axi4l_addr_t'(40'ha010_0000);

    localparam  axi4l_addr_t    ADR_CORE_ID            = axi4l_addr_t'('h00) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_CORE_VERSION       = axi4l_addr_t'('h01) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_CTL_CONTROL        = axi4l_addr_t'('h04) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_CTL_STATUS         = axi4l_addr_t'('h05) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_CTL_INDEX          = axi4l_addr_t'('h07) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_CTL_SKIP           = axi4l_addr_t'('h08) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_CTL_FRM_TIMER_EN   = axi4l_addr_t'('h0a) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_CTL_FRM_TIMEOUT    = axi4l_addr_t'('h0b) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_PARAM_WIDTH        = axi4l_addr_t'('h10) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_PARAM_HEIGHT       = axi4l_addr_t'('h11) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_PARAM_FILL         = axi4l_addr_t'('h12) * (axi4l_peri.DATA_BITS/8);
    localparam  axi4l_addr_t    ADR_PARAM_TIMEOUT      = axi4l_addr_t'('h13) * (axi4l_peri.DATA_BITS/8);

    jelly3_axi4l_accessor
            #(
                .RAND_RATE_AW   (0),
                .RAND_RATE_W    (0),
                .RAND_RATE_B    (0),
                .RAND_RATE_AR   (0),
                .RAND_RATE_R    (0)
            )
        u_axi4l_accessor
            (
                .m_axi4l        (axi4l_peri.m)
            );

    initial begin
        axi4l_data_t    rdata;
        
        #(RATE100*200);
        $display("start");
        u_axi4l_accessor.read(ADR_FMTR + ADR_CORE_ID,          rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_CORE_VERSION,     rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_CTL_CONTROL,      rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_CTL_STATUS,       rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_CTL_INDEX,        rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_CTL_SKIP,         rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_CTL_FRM_TIMER_EN, rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_CTL_FRM_TIMEOUT,  rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_PARAM_WIDTH,      rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_PARAM_HEIGHT,     rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_PARAM_FILL,       rdata);
        u_axi4l_accessor.read(ADR_FMTR + ADR_PARAM_TIMEOUT,    rdata);
                
        #(RATE100*100);
        $display("enable");
        u_axi4l_accessor.write(ADR_FMTR + ADR_PARAM_WIDTH       , SIM_IMG_WIDTH , 4'b1111);
        u_axi4l_accessor.write(ADR_FMTR + ADR_PARAM_HEIGHT      , SIM_IMG_HEIGHT, 4'b1111);
        u_axi4l_accessor.write(ADR_FMTR + ADR_PARAM_TIMEOUT     , 1000          , 4'b1111);
        u_axi4l_accessor.write(ADR_FMTR + ADR_CTL_FRM_TIMEOUT   , 100000        , 4'b1111);
        u_axi4l_accessor.write(ADR_FMTR + ADR_CTL_FRM_TIMER_EN  , 1             , 4'b1111);
        u_axi4l_accessor.write(ADR_FMTR + ADR_CTL_CONTROL       , 1             , 4'b1111);
        u_axi4l_accessor.read (ADR_FMTR + ADR_CTL_STATUS        , rdata);


    end

endmodule


`default_nettype wire


// end of file
