
`timescale 1 ns / 1 ps

module design_1
    (
        fan_en  ,
        reset_n
    );
  
  output fan_en ;
  output reset_n;

  wire fan_en;
  wire reset_n;

  assign fan_en  = 1'b0  ;

endmodule
