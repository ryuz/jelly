// ---------------------------------------------------------------------------
//  Jelly  -- the system on fpga system
//
//  Ultra96V2 udmabuf test
//
//                                 Copyright (C) 2008-2026 by Ryuji Fuchikami
//                                 https://github.com/ryuz/jelly.git
// ---------------------------------------------------------------------------

`timescale 1ns / 1ps
`default_nettype none

module hub75_driver_core
            #(
                parameter   int     CLK_DIV       = 4                           ,
                parameter   int     DISP_BITS     = 16                          ,
                parameter   type    disp_t        = logic [DISP_BITS-1:0]       ,
                parameter   int     INTERVAL_BITS = 8                           ,
                parameter   type    interval_t    = logic [INTERVAL_BITS-1:0]   ,
                parameter   int     N             = 2                           ,
                parameter   int     WIDTH         = 64                          ,
                parameter   int     HEIGHT        = 32                          ,
                parameter   int     SEL_BITS      = $clog2(HEIGHT)              ,
                parameter   type    sel_t         = logic [SEL_BITS-1:0]        ,
                parameter   int     DATA_BITS     = 8                           ,
                parameter   type    data_t        = logic [DATA_BITS-1:0]       ,
                parameter   int     SLOTS         = $bits(data_t)               ,
                parameter   int     DEPTH         = N * HEIGHT * WIDTH          ,
                parameter   int     ADDR_BITS     = $clog2(DEPTH)               ,
                parameter   type    addr_t        = logic [ADDR_BITS-1:0]       ,
                parameter           RAM_TYPE      = "block"                     ,
                parameter   bit     READMEMB      = 1'b0                        ,
                parameter   bit     READMEMH      = 1'b0                        ,
                parameter           READMEM_FILE  = ""                          
            )
            (
                input   var logic                   reset       ,
                input   var logic                   clk         ,
                input   var logic                   enable      ,
                input   var logic                   flip_h      ,
                input   var logic                   flip_v      ,
                input   var disp_t      [SLOTS-1:0] disp        ,
                input   var interval_t  [SLOTS-1:0] interval    ,

                output  var logic                   hub75_cke   ,
                output  var logic                   hub75_oe_n  ,
                output  var logic                   hub75_lat   ,
                output  var sel_t                   hub75_sel   ,
                output  var logic       [N-1:0]     hub75_r     ,
                output  var logic       [N-1:0]     hub75_g     ,
                output  var logic       [N-1:0]     hub75_b     ,

                input   var logic                   mem_clk     ,
                input   var logic                   mem_we      ,
                input   var addr_t                  mem_addr    ,
                input   var data_t                  mem_r       ,
                input   var data_t                  mem_g       ,
                input   var data_t                  mem_b       
            );
    
    localparam  int     MEM_DEPTH     = HEIGHT * WIDTH                  ;
    localparam  int     MEM_ADDR_BITS = $clog2(MEM_DEPTH)               ;
    localparam  type    mem_addr_t    = logic       [MEM_ADDR_BITS-1:0] ;
    localparam  type    mem_we_t      = logic       [N-1:0]             ;
    localparam  type    mem_word_t    = data_t      [2:0]               ;
    localparam  type    mem_data_t    = mem_word_t  [N-1:0]             ;

    mem_we_t        mem_wr_en       ;
    mem_addr_t      mem_wr_addr     ;
    mem_data_t      mem_wr_din      ;
    mem_addr_t      mem_rd_addr     ;
    mem_data_t      mem_rd_dout     ;

    jelly3_ram_simple_dualport
            #(
                .ADDR_BITS      (MEM_ADDR_BITS      ),
                .WE_BITS        (N                  ),
                .DATA_BITS      ($bits(mem_data_t)  ),
                .WORD_BITS      ($bits(mem_word_t)  ),
                .MEM_DEPTH      (MEM_DEPTH          ),
                .RAM_TYPE       (RAM_TYPE           ),
                .DOUT_REG       (1'b1               ),
                .READMEMB       (READMEMB           ),
                .READMEMH       (READMEMH           ),
                .READMEM_FILE   (READMEM_FILE       )
            )
        u_ram_simple_dualport
            (
                .wr_clk         (mem_clk            ),
                .wr_en          (mem_wr_en          ),
                .wr_addr        (mem_wr_addr        ),
                .wr_din         (mem_wr_din         ),
                
                .rd_clk         (clk                ),
                .rd_en          (1'b1               ),
                .rd_regcke      (1'b1               ),
                .rd_addr        (mem_rd_addr        ),
                .rd_dout        (mem_rd_dout        )
            );
    
    assign mem_wr_en   = mem_we ? (1 << (mem_addr >> MEM_ADDR_BITS)) : '0;
    assign mem_wr_addr = mem_addr_t'(mem_addr);
    assign mem_wr_din  = {N{mem_r, mem_g, mem_b}};

    localparam  type    div_t  = logic [$clog2(CLK_DIV)-1:0];
    localparam  type    x_t    = logic [$clog2(WIDTH )-1:0] ;
    localparam  type    y_t    = logic [$clog2(HEIGHT)-1:0] ;
    localparam  int     F_BITS = $clog2($bits(data_t))      ;
    localparam  type    f_t    = logic [F_BITS-1:0]         ;

    typedef enum {
        IDLE,
        SETUP,
        TRANS,
        LAT
    } state_t;


    // stage 0
    div_t                   st0_div     ;
    state_t                 st0_state   ;
    logic                   st0_cke     ;
    logic                   st0_lat     ;
    logic                   st0_oe_n    ;
    logic                   st0_en      ;
    sel_t                   st0_sel     ;
    x_t                     st0_x       ;
    y_t                     st0_y       ;
    f_t                     st0_f       ;
    disp_t                  st0_disp    ;
    interval_t  [SLOTS-1:0] st0_interval;

    always_ff @(posedge clk) begin
        if ( reset ) begin
            st0_div   <= '0    ;
            st0_state <= IDLE  ;
            st0_cke   <= 1'b0  ;
            st0_lat   <= 1'b0  ;
            st0_oe_n  <= 1'b1  ;
            st0_en    <= 1'b0  ;
            st0_sel   <= '0    ;
            st0_x     <= '0    ;
            st0_y     <= '0    ;
            st0_f     <= '0    ;
            st0_disp  <= '0    ;
            st0_interval <= '0  ;
        end
        else begin
            if ( st0_state == TRANS ) begin
                st0_disp <= st0_disp - 1;
                if ( st0_disp == '0 ) begin
                    st0_oe_n <= 1'b1  ;
                end
            end

            st0_div <= st0_div + 1;
            if ( st0_div == div_t'(CLK_DIV - 1) ) begin
                st0_div   <= '0     ;
                case ( st0_state )
                IDLE:
                    begin
                        if ( enable ) begin
                            st0_state <= SETUP  ;
                        end
                        st0_cke   <= 1'b0   ;
                        st0_lat   <= 1'b0   ;
                        st0_oe_n  <= 1'b1   ;
                    end
                
                SETUP:
                    begin
                        st0_state <= TRANS  ;
                        st0_cke   <= 1'b0   ;
                        st0_lat   <= 1'b0   ;
                        st0_oe_n  <= 1'b0   ;
                    end

                TRANS:
                    begin
                        st0_cke <= ~st0_cke;
                        if ( st0_cke ) begin
                            st0_x <= st0_x + 1;
                            if ( st0_x == x_t'(WIDTH-1) ) begin
                                st0_state <= LAT    ;
                                st0_lat   <= 1'b1   ;
                                st0_oe_n  <= 1'b1   ;
                                st0_sel   <= st0_y  ;
                                st0_x     <= '0     ;
                                st0_y     <= st0_y + 1;
                                st0_disp  <= disp[st0_f];
                                if ( st0_interval[st0_f] == 0 ) begin
                                    st0_en <= 1'b1;
                                end
                                else begin
                                    st0_en <= 1'b0;
                                end
                                if ( st0_y == y_t'(HEIGHT-1) ) begin
                                    st0_y   <= '0;
                                    st0_f   <= st0_f + 1;
                                    if ( st0_f == f_t'($bits(data_t)-1) ) begin
                                        st0_f <= '0;
                                        for ( int i = 0; i < SLOTS; i++ ) begin
                                            st0_interval[i] <= st0_interval[i] - 1;
                                            if ( st0_interval[i] == 0 ) begin
                                                st0_interval[i] <= interval[i];
                                            end
                                        end
                                    end
                                end
                            end
                        end
                    end

                LAT:
                    begin
                        st0_state <= IDLE   ;
                        st0_lat   <= 1'b1   ;
                        st0_oe_n  <= 1'b1   ;
                    end
                endcase
            end
        end
    end

    x_t         mem_x       ;
    y_t         mem_y       ;
    assign mem_x = flip_h ? ~st0_x : st0_x;
    assign mem_y = flip_v ? ~st0_y : st0_y;
    assign mem_rd_addr = {mem_y, mem_x};

    logic           st1_cke ;
    logic           st1_lat ;
    logic           st1_oe_n;
    sel_t           st1_sel ;
    f_t             st1_f   ;

    logic           st2_cke ;
    logic           st2_lat ;
    logic           st2_oe_n;
    sel_t           st2_sel ;
    f_t             st2_f   ;

    logic           st3_cke ;
    logic           st3_lat ;
    logic           st3_oe_n;
    sel_t           st3_sel ;
    logic   [N-1:0] st3_r   ;
    logic   [N-1:0] st3_g   ;
    logic   [N-1:0] st3_b   ;

    always_ff @(posedge clk) begin
        st1_cke  <= st0_cke ;
        st1_lat  <= st0_lat ;
        st1_oe_n <= st0_oe_n | ~st0_en;
        st1_sel  <= st0_sel ;
        st1_f    <= st0_f   ;

        st2_cke  <= st1_cke ;
        st2_lat  <= st1_lat ;
        st2_oe_n <= st1_oe_n;
        st2_sel  <= st1_sel ;
        st2_f    <= st1_f   ;

        st3_cke  <= st2_cke ;
        st3_lat  <= st2_lat ;
        st3_oe_n <= st2_oe_n;
        st3_sel  <= st2_sel ;
        st3_r    <= '0;
        st3_g    <= '0;
        st3_b    <= '0;
//      if ( st2_f >= 0 ) begin
            for ( int i = 0; i < N; i++ ) begin
                st3_r[i] <= mem_rd_dout[i][2][st2_f];
                st3_g[i] <= mem_rd_dout[i][1][st2_f];
                st3_b[i] <= mem_rd_dout[i][0][st2_f];
            end
//      end
    end

    assign  hub75_cke  = st3_cke ;
    assign  hub75_oe_n = st3_oe_n;
    assign  hub75_lat  = st3_lat ;
    assign  hub75_sel  = st3_sel ;
    assign  hub75_r    = st3_r   ;
    assign  hub75_g    = st3_g   ;
    assign  hub75_b    = st3_b   ;

endmodule



`default_nettype wire


// end of file
