// ---------------------------------------------------------------------------
//  Jelly  -- the system on fpga system
//
//  Test DMA
//
//                                 Copyright (C) 2008-2020 by Ryuji Fuchikami
//                                 https://github.com/ryuz/jelly.git
// ---------------------------------------------------------------------------


`timescale 1ns / 1ps
`default_nettype none


module sin_3phase_tbl
        (
            input   wire            reset,
            input   wire            clk,
            input   wire            cke,
            
            input   wire    [9:0]   in_phase,
            
            output  wire    [11:0]  out_x,
            output  wire    [11:0]  out_y,
            output  wire    [11:0]  out_z
        );
    
    reg     [35:0]  dout;
    always @(posedge clk) begin
        if ( cke ) begin
            case ( in_phase )
            10'd0000: dout <= 36'b000100010011_111011101101_100000000000;
            10'd0001: dout <= 36'b000100001101_111011100110_100000001101;
            10'd0002: dout <= 36'b000100000111_111011100000_100000011001;
            10'd0003: dout <= 36'b000100000001_111011011010_100000100110;
            10'd0004: dout <= 36'b000011111011_111011010011_100000110010;
            10'd0005: dout <= 36'b000011110101_111011001101_100000111111;
            10'd0006: dout <= 36'b000011101111_111011000110_100001001011;
            10'd0007: dout <= 36'b000011101001_111010111111_100001011000;
            10'd0008: dout <= 36'b000011100011_111010111000_100001100100;
            10'd0009: dout <= 36'b000011011101_111010110010_100001110001;
            10'd0010: dout <= 36'b000011011000_111010101011_100001111110;
            10'd0011: dout <= 36'b000011010010_111010100100_100010001010;
            10'd0012: dout <= 36'b000011001101_111010011101_100010010111;
            10'd0013: dout <= 36'b000011000111_111010010110_100010100011;
            10'd0014: dout <= 36'b000011000010_111010001110_100010110000;
            10'd0015: dout <= 36'b000010111101_111010000111_100010111100;
            10'd0016: dout <= 36'b000010110111_111010000000_100011001001;
            10'd0017: dout <= 36'b000010110010_111001111001_100011010101;
            10'd0018: dout <= 36'b000010101101_111001110001_100011100010;
            10'd0019: dout <= 36'b000010101000_111001101010_100011101110;
            10'd0020: dout <= 36'b000010100011_111001100010_100011111011;
            10'd0021: dout <= 36'b000010011110_111001011011_100100000111;
            10'd0022: dout <= 36'b000010011010_111001010011_100100010011;
            10'd0023: dout <= 36'b000010010101_111001001011_100100100000;
            10'd0024: dout <= 36'b000010010000_111001000011_100100101100;
            10'd0025: dout <= 36'b000010001100_111000111100_100100111001;
            10'd0026: dout <= 36'b000010000111_111000110100_100101000101;
            10'd0027: dout <= 36'b000010000011_111000101100_100101010010;
            10'd0028: dout <= 36'b000001111110_111000100100_100101011110;
            10'd0029: dout <= 36'b000001111010_111000011100_100101101010;
            10'd0030: dout <= 36'b000001110110_111000010011_100101110111;
            10'd0031: dout <= 36'b000001110010_111000001011_100110000011;
            10'd0032: dout <= 36'b000001101110_111000000011_100110001111;
            10'd0033: dout <= 36'b000001101010_110111111011_100110011100;
            10'd0034: dout <= 36'b000001100110_110111110010_100110101000;
            10'd0035: dout <= 36'b000001100010_110111101010_100110110100;
            10'd0036: dout <= 36'b000001011110_110111100001_100111000001;
            10'd0037: dout <= 36'b000001011010_110111011001_100111001101;
            10'd0038: dout <= 36'b000001010111_110111010000_100111011001;
            10'd0039: dout <= 36'b000001010011_110111001000_100111100101;
            10'd0040: dout <= 36'b000001010000_110110111111_100111110001;
            10'd0041: dout <= 36'b000001001100_110110110110_100111111110;
            10'd0042: dout <= 36'b000001001001_110110101101_101000001010;
            10'd0043: dout <= 36'b000001000110_110110100100_101000010110;
            10'd0044: dout <= 36'b000001000010_110110011100_101000100010;
            10'd0045: dout <= 36'b000000111111_110110010011_101000101110;
            10'd0046: dout <= 36'b000000111100_110110001010_101000111010;
            10'd0047: dout <= 36'b000000111001_110110000000_101001000110;
            10'd0048: dout <= 36'b000000110110_110101110111_101001010010;
            10'd0049: dout <= 36'b000000110100_110101101110_101001011110;
            10'd0050: dout <= 36'b000000110001_110101100101_101001101010;
            10'd0051: dout <= 36'b000000101110_110101011100_101001110110;
            10'd0052: dout <= 36'b000000101100_110101010010_101010000010;
            10'd0053: dout <= 36'b000000101001_110101001001_101010001110;
            10'd0054: dout <= 36'b000000100111_110100111111_101010011010;
            10'd0055: dout <= 36'b000000100100_110100110110_101010100110;
            10'd0056: dout <= 36'b000000100010_110100101100_101010110010;
            10'd0057: dout <= 36'b000000100000_110100100011_101010111101;
            10'd0058: dout <= 36'b000000011110_110100011001_101011001001;
            10'd0059: dout <= 36'b000000011100_110100001111_101011010101;
            10'd0060: dout <= 36'b000000011010_110100000110_101011100001;
            10'd0061: dout <= 36'b000000011000_110011111100_101011101100;
            10'd0062: dout <= 36'b000000010110_110011110010_101011111000;
            10'd0063: dout <= 36'b000000010100_110011101000_101100000100;
            10'd0064: dout <= 36'b000000010011_110011011110_101100001111;
            10'd0065: dout <= 36'b000000010001_110011010100_101100011011;
            10'd0066: dout <= 36'b000000001111_110011001010_101100100111;
            10'd0067: dout <= 36'b000000001110_110011000000_101100110010;
            10'd0068: dout <= 36'b000000001101_110010110110_101100111110;
            10'd0069: dout <= 36'b000000001011_110010101100_101101001001;
            10'd0070: dout <= 36'b000000001010_110010100010_101101010100;
            10'd0071: dout <= 36'b000000001001_110010010111_101101100000;
            10'd0072: dout <= 36'b000000001000_110010001101_101101101011;
            10'd0073: dout <= 36'b000000000111_110010000011_101101110111;
            10'd0074: dout <= 36'b000000000110_110001111000_101110000010;
            10'd0075: dout <= 36'b000000000101_110001101110_101110001101;
            10'd0076: dout <= 36'b000000000100_110001100011_101110011000;
            10'd0077: dout <= 36'b000000000100_110001011001_101110100100;
            10'd0078: dout <= 36'b000000000011_110001001110_101110101111;
            10'd0079: dout <= 36'b000000000011_110001000100_101110111010;
            10'd0080: dout <= 36'b000000000010_110000111001_101111000101;
            10'd0081: dout <= 36'b000000000010_110000101110_101111010000;
            10'd0082: dout <= 36'b000000000001_110000100100_101111011011;
            10'd0083: dout <= 36'b000000000001_110000011001_101111100110;
            10'd0084: dout <= 36'b000000000001_110000001110_101111110001;
            10'd0085: dout <= 36'b000000000001_110000000011_101111111100;
            10'd0086: dout <= 36'b000000000001_101111111000_110000000111;
            10'd0087: dout <= 36'b000000000001_101111101101_110000010010;
            10'd0088: dout <= 36'b000000000001_101111100010_110000011100;
            10'd0089: dout <= 36'b000000000010_101111010111_110000100111;
            10'd0090: dout <= 36'b000000000010_101111001100_110000110010;
            10'd0091: dout <= 36'b000000000010_101111000001_110000111101;
            10'd0092: dout <= 36'b000000000011_101110110110_110001000111;
            10'd0093: dout <= 36'b000000000011_101110101011_110001010010;
            10'd0094: dout <= 36'b000000000100_101110100000_110001011100;
            10'd0095: dout <= 36'b000000000101_101110010101_110001100111;
            10'd0096: dout <= 36'b000000000101_101110001001_110001110001;
            10'd0097: dout <= 36'b000000000110_101101111110_110001111100;
            10'd0098: dout <= 36'b000000000111_101101110011_110010000110;
            10'd0099: dout <= 36'b000000001000_101101100111_110010010000;
            10'd0100: dout <= 36'b000000001001_101101011100_110010011011;
            10'd0101: dout <= 36'b000000001010_101101010001_110010100101;
            10'd0102: dout <= 36'b000000001100_101101000101_110010101111;
            10'd0103: dout <= 36'b000000001101_101100111010_110010111001;
            10'd0104: dout <= 36'b000000001110_101100101110_110011000011;
            10'd0105: dout <= 36'b000000010000_101100100011_110011001101;
            10'd0106: dout <= 36'b000000010001_101100010111_110011010111;
            10'd0107: dout <= 36'b000000010011_101100001011_110011100001;
            10'd0108: dout <= 36'b000000010101_101100000000_110011101011;
            10'd0109: dout <= 36'b000000010111_101011110100_110011110101;
            10'd0110: dout <= 36'b000000011000_101011101001_110011111111;
            10'd0111: dout <= 36'b000000011010_101011011101_110100001001;
            10'd0112: dout <= 36'b000000011100_101011010001_110100010011;
            10'd0113: dout <= 36'b000000011110_101011000101_110100011100;
            10'd0114: dout <= 36'b000000100001_101010111001_110100100110;
            10'd0115: dout <= 36'b000000100011_101010101110_110100110000;
            10'd0116: dout <= 36'b000000100101_101010100010_110100111001;
            10'd0117: dout <= 36'b000000101000_101010010110_110101000011;
            10'd0118: dout <= 36'b000000101010_101010001010_110101001100;
            10'd0119: dout <= 36'b000000101101_101001111110_110101010101;
            10'd0120: dout <= 36'b000000101111_101001110010_110101011111;
            10'd0121: dout <= 36'b000000110010_101001100110_110101101000;
            10'd0122: dout <= 36'b000000110101_101001011010_110101110001;
            10'd0123: dout <= 36'b000000110111_101001001110_110101111010;
            10'd0124: dout <= 36'b000000111010_101001000010_110110000011;
            10'd0125: dout <= 36'b000000111101_101000110110_110110001101;
            10'd0126: dout <= 36'b000001000000_101000101010_110110010110;
            10'd0127: dout <= 36'b000001000100_101000011110_110110011111;
            10'd0128: dout <= 36'b000001000111_101000010010_110110100111;
            10'd0129: dout <= 36'b000001001010_101000000110_110110110000;
            10'd0130: dout <= 36'b000001001101_100111111001_110110111001;
            10'd0131: dout <= 36'b000001010001_100111101101_110111000010;
            10'd0132: dout <= 36'b000001010100_100111100001_110111001011;
            10'd0133: dout <= 36'b000001011000_100111010101_110111010011;
            10'd0134: dout <= 36'b000001011100_100111001001_110111011100;
            10'd0135: dout <= 36'b000001011111_100110111100_110111100100;
            10'd0136: dout <= 36'b000001100011_100110110000_110111101101;
            10'd0137: dout <= 36'b000001100111_100110100100_110111110101;
            10'd0138: dout <= 36'b000001101011_100110011000_110111111101;
            10'd0139: dout <= 36'b000001101111_100110001011_111000000110;
            10'd0140: dout <= 36'b000001110011_100101111111_111000001110;
            10'd0141: dout <= 36'b000001110111_100101110011_111000010110;
            10'd0142: dout <= 36'b000001111011_100101100110_111000011110;
            10'd0143: dout <= 36'b000010000000_100101011010_111000100110;
            10'd0144: dout <= 36'b000010000100_100101001101_111000101110;
            10'd0145: dout <= 36'b000010001001_100101000001_111000110110;
            10'd0146: dout <= 36'b000010001101_100100110101_111000111110;
            10'd0147: dout <= 36'b000010010010_100100101000_111001000110;
            10'd0148: dout <= 36'b000010010110_100100011100_111001001110;
            10'd0149: dout <= 36'b000010011011_100100001111_111001010101;
            10'd0150: dout <= 36'b000010100000_100100000011_111001011101;
            10'd0151: dout <= 36'b000010100101_100011110110_111001100101;
            10'd0152: dout <= 36'b000010101010_100011101010_111001101100;
            10'd0153: dout <= 36'b000010101111_100011011101_111001110100;
            10'd0154: dout <= 36'b000010110100_100011010001_111001111011;
            10'd0155: dout <= 36'b000010111001_100011000100_111010000010;
            10'd0156: dout <= 36'b000010111110_100010111000_111010001010;
            10'd0157: dout <= 36'b000011000100_100010101011_111010010001;
            10'd0158: dout <= 36'b000011001001_100010011111_111010011000;
            10'd0159: dout <= 36'b000011001111_100010010010_111010011111;
            10'd0160: dout <= 36'b000011010100_100010000110_111010100110;
            10'd0161: dout <= 36'b000011011010_100001111001_111010101101;
            10'd0162: dout <= 36'b000011011111_100001101101_111010110100;
            10'd0163: dout <= 36'b000011100101_100001100000_111010111011;
            10'd0164: dout <= 36'b000011101011_100001010100_111011000001;
            10'd0165: dout <= 36'b000011110001_100001000111_111011001000;
            10'd0166: dout <= 36'b000011110111_100000111011_111011001111;
            10'd0167: dout <= 36'b000011111101_100000101110_111011010101;
            10'd0168: dout <= 36'b000100000011_100000100001_111011011100;
            10'd0169: dout <= 36'b000100001001_100000010101_111011100010;
            10'd0170: dout <= 36'b000100001111_100000001000_111011101001;
            10'd0171: dout <= 36'b000100010101_011111111100_111011101111;
            10'd0172: dout <= 36'b000100011100_011111101111_111011110101;
            10'd0173: dout <= 36'b000100100010_011111100011_111011111011;
            10'd0174: dout <= 36'b000100101001_011111010110_111100000001;
            10'd0175: dout <= 36'b000100101111_011111001010_111100000111;
            10'd0176: dout <= 36'b000100110110_011110111101_111100001101;
            10'd0177: dout <= 36'b000100111100_011110110000_111100010011;
            10'd0178: dout <= 36'b000101000011_011110100100_111100011001;
            10'd0179: dout <= 36'b000101001010_011110010111_111100011111;
            10'd0180: dout <= 36'b000101010001_011110001011_111100100100;
            10'd0181: dout <= 36'b000101011000_011101111110_111100101010;
            10'd0182: dout <= 36'b000101011111_011101110010_111100110000;
            10'd0183: dout <= 36'b000101100110_011101100101_111100110101;
            10'd0184: dout <= 36'b000101101101_011101011001_111100111010;
            10'd0185: dout <= 36'b000101110100_011101001100_111101000000;
            10'd0186: dout <= 36'b000101111011_011101000000_111101000101;
            10'd0187: dout <= 36'b000110000011_011100110011_111101001010;
            10'd0188: dout <= 36'b000110001010_011100100111_111101001111;
            10'd0189: dout <= 36'b000110010001_011100011010_111101010100;
            10'd0190: dout <= 36'b000110011001_011100001110_111101011001;
            10'd0191: dout <= 36'b000110100000_011100000001_111101011110;
            10'd0192: dout <= 36'b000110101000_011011110101_111101100011;
            10'd0193: dout <= 36'b000110110000_011011101000_111101101000;
            10'd0194: dout <= 36'b000110110111_011011011100_111101101101;
            10'd0195: dout <= 36'b000110111111_011011010000_111101110001;
            10'd0196: dout <= 36'b000111000111_011011000011_111101110110;
            10'd0197: dout <= 36'b000111001111_011010110111_111101111010;
            10'd0198: dout <= 36'b000111010111_011010101010_111101111111;
            10'd0199: dout <= 36'b000111011111_011010011110_111110000011;
            10'd0200: dout <= 36'b000111100111_011010010010_111110000111;
            10'd0201: dout <= 36'b000111101111_011010000101_111110001100;
            10'd0202: dout <= 36'b000111110111_011001111001_111110010000;
            10'd0203: dout <= 36'b001000000000_011001101101_111110010100;
            10'd0204: dout <= 36'b001000001000_011001100000_111110011000;
            10'd0205: dout <= 36'b001000010000_011001010100_111110011100;
            10'd0206: dout <= 36'b001000011001_011001001000_111110011111;
            10'd0207: dout <= 36'b001000100001_011000111011_111110100011;
            10'd0208: dout <= 36'b001000101010_011000101111_111110100111;
            10'd0209: dout <= 36'b001000110011_011000100011_111110101010;
            10'd0210: dout <= 36'b001000111011_011000010111_111110101110;
            10'd0211: dout <= 36'b001001000100_011000001011_111110110001;
            10'd0212: dout <= 36'b001001001101_010111111110_111110110101;
            10'd0213: dout <= 36'b001001010110_010111110010_111110111000;
            10'd0214: dout <= 36'b001001011110_010111100110_111110111011;
            10'd0215: dout <= 36'b001001100111_010111011010_111110111111;
            10'd0216: dout <= 36'b001001110000_010111001110_111111000010;
            10'd0217: dout <= 36'b001001111001_010111000010_111111000101;
            10'd0218: dout <= 36'b001010000011_010110110110_111111001000;
            10'd0219: dout <= 36'b001010001100_010110101010_111111001010;
            10'd0220: dout <= 36'b001010010101_010110011110_111111001101;
            10'd0221: dout <= 36'b001010011110_010110010010_111111010000;
            10'd0222: dout <= 36'b001010101000_010110000110_111111010011;
            10'd0223: dout <= 36'b001010110001_010101111010_111111010101;
            10'd0224: dout <= 36'b001010111010_010101101110_111111011000;
            10'd0225: dout <= 36'b001011000100_010101100010_111111011010;
            10'd0226: dout <= 36'b001011001101_010101010110_111111011100;
            10'd0227: dout <= 36'b001011010111_010101001010_111111011111;
            10'd0228: dout <= 36'b001011100000_010100111111_111111100001;
            10'd0229: dout <= 36'b001011101010_010100110011_111111100011;
            10'd0230: dout <= 36'b001011110100_010100100111_111111100101;
            10'd0231: dout <= 36'b001011111110_010100011011_111111100111;
            10'd0232: dout <= 36'b001100000111_010100010000_111111101001;
            10'd0233: dout <= 36'b001100010001_010100000100_111111101011;
            10'd0234: dout <= 36'b001100011011_010011111000_111111101100;
            10'd0235: dout <= 36'b001100100101_010011101101_111111101110;
            10'd0236: dout <= 36'b001100101111_010011100001_111111110000;
            10'd0237: dout <= 36'b001100111001_010011010110_111111110001;
            10'd0238: dout <= 36'b001101000011_010011001010_111111110011;
            10'd0239: dout <= 36'b001101001101_010010111111_111111110100;
            10'd0240: dout <= 36'b001101011000_010010110011_111111110101;
            10'd0241: dout <= 36'b001101100010_010010101000_111111110110;
            10'd0242: dout <= 36'b001101101100_010010011100_111111110111;
            10'd0243: dout <= 36'b001101110110_010010010001_111111111000;
            10'd0244: dout <= 36'b001110000001_010010000110_111111111001;
            10'd0245: dout <= 36'b001110001011_010001111010_111111111010;
            10'd0246: dout <= 36'b001110010110_010001101111_111111111011;
            10'd0247: dout <= 36'b001110100000_010001100100_111111111100;
            10'd0248: dout <= 36'b001110101011_010001011001_111111111101;
            10'd0249: dout <= 36'b001110110101_010001001110_111111111101;
            10'd0250: dout <= 36'b001111000000_010001000010_111111111110;
            10'd0251: dout <= 36'b001111001011_010000110111_111111111110;
            10'd0252: dout <= 36'b001111010101_010000101100_111111111110;
            10'd0253: dout <= 36'b001111100000_010000100001_111111111111;
            10'd0254: dout <= 36'b001111101011_010000010110_111111111111;
            10'd0255: dout <= 36'b001111110110_010000001011_111111111111;
            10'd0256: dout <= 36'b010000000000_010000000001_111111111111;
            10'd0257: dout <= 36'b010000001011_001111110110_111111111111;
            10'd0258: dout <= 36'b010000010110_001111101011_111111111111;
            10'd0259: dout <= 36'b010000100001_001111100000_111111111111;
            10'd0260: dout <= 36'b010000101100_001111010101_111111111110;
            10'd0261: dout <= 36'b010000110111_001111001011_111111111110;
            10'd0262: dout <= 36'b010001000010_001111000000_111111111110;
            10'd0263: dout <= 36'b010001001110_001110110101_111111111101;
            10'd0264: dout <= 36'b010001011001_001110101011_111111111101;
            10'd0265: dout <= 36'b010001100100_001110100000_111111111100;
            10'd0266: dout <= 36'b010001101111_001110010110_111111111011;
            10'd0267: dout <= 36'b010001111010_001110001011_111111111010;
            10'd0268: dout <= 36'b010010000110_001110000001_111111111001;
            10'd0269: dout <= 36'b010010010001_001101110110_111111111000;
            10'd0270: dout <= 36'b010010011100_001101101100_111111110111;
            10'd0271: dout <= 36'b010010101000_001101100010_111111110110;
            10'd0272: dout <= 36'b010010110011_001101011000_111111110101;
            10'd0273: dout <= 36'b010010111111_001101001101_111111110100;
            10'd0274: dout <= 36'b010011001010_001101000011_111111110011;
            10'd0275: dout <= 36'b010011010110_001100111001_111111110001;
            10'd0276: dout <= 36'b010011100001_001100101111_111111110000;
            10'd0277: dout <= 36'b010011101101_001100100101_111111101110;
            10'd0278: dout <= 36'b010011111000_001100011011_111111101100;
            10'd0279: dout <= 36'b010100000100_001100010001_111111101011;
            10'd0280: dout <= 36'b010100010000_001100000111_111111101001;
            10'd0281: dout <= 36'b010100011011_001011111110_111111100111;
            10'd0282: dout <= 36'b010100100111_001011110100_111111100101;
            10'd0283: dout <= 36'b010100110011_001011101010_111111100011;
            10'd0284: dout <= 36'b010100111111_001011100000_111111100001;
            10'd0285: dout <= 36'b010101001010_001011010111_111111011111;
            10'd0286: dout <= 36'b010101010110_001011001101_111111011100;
            10'd0287: dout <= 36'b010101100010_001011000100_111111011010;
            10'd0288: dout <= 36'b010101101110_001010111010_111111011000;
            10'd0289: dout <= 36'b010101111010_001010110001_111111010101;
            10'd0290: dout <= 36'b010110000110_001010101000_111111010011;
            10'd0291: dout <= 36'b010110010010_001010011110_111111010000;
            10'd0292: dout <= 36'b010110011110_001010010101_111111001101;
            10'd0293: dout <= 36'b010110101010_001010001100_111111001010;
            10'd0294: dout <= 36'b010110110110_001010000011_111111001000;
            10'd0295: dout <= 36'b010111000010_001001111001_111111000101;
            10'd0296: dout <= 36'b010111001110_001001110000_111111000010;
            10'd0297: dout <= 36'b010111011010_001001100111_111110111111;
            10'd0298: dout <= 36'b010111100110_001001011110_111110111011;
            10'd0299: dout <= 36'b010111110010_001001010110_111110111000;
            10'd0300: dout <= 36'b010111111110_001001001101_111110110101;
            10'd0301: dout <= 36'b011000001011_001001000100_111110110001;
            10'd0302: dout <= 36'b011000010111_001000111011_111110101110;
            10'd0303: dout <= 36'b011000100011_001000110011_111110101010;
            10'd0304: dout <= 36'b011000101111_001000101010_111110100111;
            10'd0305: dout <= 36'b011000111011_001000100001_111110100011;
            10'd0306: dout <= 36'b011001001000_001000011001_111110011111;
            10'd0307: dout <= 36'b011001010100_001000010000_111110011100;
            10'd0308: dout <= 36'b011001100000_001000001000_111110011000;
            10'd0309: dout <= 36'b011001101101_001000000000_111110010100;
            10'd0310: dout <= 36'b011001111001_000111110111_111110010000;
            10'd0311: dout <= 36'b011010000101_000111101111_111110001100;
            10'd0312: dout <= 36'b011010010010_000111100111_111110000111;
            10'd0313: dout <= 36'b011010011110_000111011111_111110000011;
            10'd0314: dout <= 36'b011010101010_000111010111_111101111111;
            10'd0315: dout <= 36'b011010110111_000111001111_111101111010;
            10'd0316: dout <= 36'b011011000011_000111000111_111101110110;
            10'd0317: dout <= 36'b011011010000_000110111111_111101110001;
            10'd0318: dout <= 36'b011011011100_000110110111_111101101101;
            10'd0319: dout <= 36'b011011101000_000110110000_111101101000;
            10'd0320: dout <= 36'b011011110101_000110101000_111101100011;
            10'd0321: dout <= 36'b011100000001_000110100000_111101011110;
            10'd0322: dout <= 36'b011100001110_000110011001_111101011001;
            10'd0323: dout <= 36'b011100011010_000110010001_111101010100;
            10'd0324: dout <= 36'b011100100111_000110001010_111101001111;
            10'd0325: dout <= 36'b011100110011_000110000011_111101001010;
            10'd0326: dout <= 36'b011101000000_000101111011_111101000101;
            10'd0327: dout <= 36'b011101001100_000101110100_111101000000;
            10'd0328: dout <= 36'b011101011001_000101101101_111100111010;
            10'd0329: dout <= 36'b011101100101_000101100110_111100110101;
            10'd0330: dout <= 36'b011101110010_000101011111_111100110000;
            10'd0331: dout <= 36'b011101111110_000101011000_111100101010;
            10'd0332: dout <= 36'b011110001011_000101010001_111100100100;
            10'd0333: dout <= 36'b011110010111_000101001010_111100011111;
            10'd0334: dout <= 36'b011110100100_000101000011_111100011001;
            10'd0335: dout <= 36'b011110110000_000100111100_111100010011;
            10'd0336: dout <= 36'b011110111101_000100110110_111100001101;
            10'd0337: dout <= 36'b011111001010_000100101111_111100000111;
            10'd0338: dout <= 36'b011111010110_000100101001_111100000001;
            10'd0339: dout <= 36'b011111100011_000100100010_111011111011;
            10'd0340: dout <= 36'b011111101111_000100011100_111011110101;
            10'd0341: dout <= 36'b011111111100_000100010101_111011101111;
            10'd0342: dout <= 36'b100000001000_000100001111_111011101001;
            10'd0343: dout <= 36'b100000010101_000100001001_111011100010;
            10'd0344: dout <= 36'b100000100001_000100000011_111011011100;
            10'd0345: dout <= 36'b100000101110_000011111101_111011010101;
            10'd0346: dout <= 36'b100000111011_000011110111_111011001111;
            10'd0347: dout <= 36'b100001000111_000011110001_111011001000;
            10'd0348: dout <= 36'b100001010100_000011101011_111011000001;
            10'd0349: dout <= 36'b100001100000_000011100101_111010111011;
            10'd0350: dout <= 36'b100001101101_000011011111_111010110100;
            10'd0351: dout <= 36'b100001111001_000011011010_111010101101;
            10'd0352: dout <= 36'b100010000110_000011010100_111010100110;
            10'd0353: dout <= 36'b100010010010_000011001111_111010011111;
            10'd0354: dout <= 36'b100010011111_000011001001_111010011000;
            10'd0355: dout <= 36'b100010101011_000011000100_111010010001;
            10'd0356: dout <= 36'b100010111000_000010111110_111010001010;
            10'd0357: dout <= 36'b100011000100_000010111001_111010000010;
            10'd0358: dout <= 36'b100011010001_000010110100_111001111011;
            10'd0359: dout <= 36'b100011011101_000010101111_111001110100;
            10'd0360: dout <= 36'b100011101010_000010101010_111001101100;
            10'd0361: dout <= 36'b100011110110_000010100101_111001100101;
            10'd0362: dout <= 36'b100100000011_000010100000_111001011101;
            10'd0363: dout <= 36'b100100001111_000010011011_111001010101;
            10'd0364: dout <= 36'b100100011100_000010010110_111001001110;
            10'd0365: dout <= 36'b100100101000_000010010010_111001000110;
            10'd0366: dout <= 36'b100100110101_000010001101_111000111110;
            10'd0367: dout <= 36'b100101000001_000010001001_111000110110;
            10'd0368: dout <= 36'b100101001101_000010000100_111000101110;
            10'd0369: dout <= 36'b100101011010_000010000000_111000100110;
            10'd0370: dout <= 36'b100101100110_000001111011_111000011110;
            10'd0371: dout <= 36'b100101110011_000001110111_111000010110;
            10'd0372: dout <= 36'b100101111111_000001110011_111000001110;
            10'd0373: dout <= 36'b100110001011_000001101111_111000000110;
            10'd0374: dout <= 36'b100110011000_000001101011_110111111101;
            10'd0375: dout <= 36'b100110100100_000001100111_110111110101;
            10'd0376: dout <= 36'b100110110000_000001100011_110111101101;
            10'd0377: dout <= 36'b100110111100_000001011111_110111100100;
            10'd0378: dout <= 36'b100111001001_000001011100_110111011100;
            10'd0379: dout <= 36'b100111010101_000001011000_110111010011;
            10'd0380: dout <= 36'b100111100001_000001010100_110111001011;
            10'd0381: dout <= 36'b100111101101_000001010001_110111000010;
            10'd0382: dout <= 36'b100111111001_000001001101_110110111001;
            10'd0383: dout <= 36'b101000000110_000001001010_110110110000;
            10'd0384: dout <= 36'b101000010010_000001000111_110110100111;
            10'd0385: dout <= 36'b101000011110_000001000100_110110011111;
            10'd0386: dout <= 36'b101000101010_000001000000_110110010110;
            10'd0387: dout <= 36'b101000110110_000000111101_110110001101;
            10'd0388: dout <= 36'b101001000010_000000111010_110110000011;
            10'd0389: dout <= 36'b101001001110_000000110111_110101111010;
            10'd0390: dout <= 36'b101001011010_000000110101_110101110001;
            10'd0391: dout <= 36'b101001100110_000000110010_110101101000;
            10'd0392: dout <= 36'b101001110010_000000101111_110101011111;
            10'd0393: dout <= 36'b101001111110_000000101101_110101010101;
            10'd0394: dout <= 36'b101010001010_000000101010_110101001100;
            10'd0395: dout <= 36'b101010010110_000000101000_110101000011;
            10'd0396: dout <= 36'b101010100010_000000100101_110100111001;
            10'd0397: dout <= 36'b101010101110_000000100011_110100110000;
            10'd0398: dout <= 36'b101010111001_000000100001_110100100110;
            10'd0399: dout <= 36'b101011000101_000000011110_110100011100;
            10'd0400: dout <= 36'b101011010001_000000011100_110100010011;
            10'd0401: dout <= 36'b101011011101_000000011010_110100001001;
            10'd0402: dout <= 36'b101011101001_000000011000_110011111111;
            10'd0403: dout <= 36'b101011110100_000000010111_110011110101;
            10'd0404: dout <= 36'b101100000000_000000010101_110011101011;
            10'd0405: dout <= 36'b101100001011_000000010011_110011100001;
            10'd0406: dout <= 36'b101100010111_000000010001_110011010111;
            10'd0407: dout <= 36'b101100100011_000000010000_110011001101;
            10'd0408: dout <= 36'b101100101110_000000001110_110011000011;
            10'd0409: dout <= 36'b101100111010_000000001101_110010111001;
            10'd0410: dout <= 36'b101101000101_000000001100_110010101111;
            10'd0411: dout <= 36'b101101010001_000000001010_110010100101;
            10'd0412: dout <= 36'b101101011100_000000001001_110010011011;
            10'd0413: dout <= 36'b101101100111_000000001000_110010010000;
            10'd0414: dout <= 36'b101101110011_000000000111_110010000110;
            10'd0415: dout <= 36'b101101111110_000000000110_110001111100;
            10'd0416: dout <= 36'b101110001001_000000000101_110001110001;
            10'd0417: dout <= 36'b101110010101_000000000101_110001100111;
            10'd0418: dout <= 36'b101110100000_000000000100_110001011100;
            10'd0419: dout <= 36'b101110101011_000000000011_110001010010;
            10'd0420: dout <= 36'b101110110110_000000000011_110001000111;
            10'd0421: dout <= 36'b101111000001_000000000010_110000111101;
            10'd0422: dout <= 36'b101111001100_000000000010_110000110010;
            10'd0423: dout <= 36'b101111010111_000000000010_110000100111;
            10'd0424: dout <= 36'b101111100010_000000000001_110000011100;
            10'd0425: dout <= 36'b101111101101_000000000001_110000010010;
            10'd0426: dout <= 36'b101111111000_000000000001_110000000111;
            10'd0427: dout <= 36'b110000000011_000000000001_101111111100;
            10'd0428: dout <= 36'b110000001110_000000000001_101111110001;
            10'd0429: dout <= 36'b110000011001_000000000001_101111100110;
            10'd0430: dout <= 36'b110000100100_000000000001_101111011011;
            10'd0431: dout <= 36'b110000101110_000000000010_101111010000;
            10'd0432: dout <= 36'b110000111001_000000000010_101111000101;
            10'd0433: dout <= 36'b110001000100_000000000011_101110111010;
            10'd0434: dout <= 36'b110001001110_000000000011_101110101111;
            10'd0435: dout <= 36'b110001011001_000000000100_101110100100;
            10'd0436: dout <= 36'b110001100011_000000000100_101110011000;
            10'd0437: dout <= 36'b110001101110_000000000101_101110001101;
            10'd0438: dout <= 36'b110001111000_000000000110_101110000010;
            10'd0439: dout <= 36'b110010000011_000000000111_101101110111;
            10'd0440: dout <= 36'b110010001101_000000001000_101101101011;
            10'd0441: dout <= 36'b110010010111_000000001001_101101100000;
            10'd0442: dout <= 36'b110010100010_000000001010_101101010100;
            10'd0443: dout <= 36'b110010101100_000000001011_101101001001;
            10'd0444: dout <= 36'b110010110110_000000001101_101100111110;
            10'd0445: dout <= 36'b110011000000_000000001110_101100110010;
            10'd0446: dout <= 36'b110011001010_000000001111_101100100111;
            10'd0447: dout <= 36'b110011010100_000000010001_101100011011;
            10'd0448: dout <= 36'b110011011110_000000010011_101100001111;
            10'd0449: dout <= 36'b110011101000_000000010100_101100000100;
            10'd0450: dout <= 36'b110011110010_000000010110_101011111000;
            10'd0451: dout <= 36'b110011111100_000000011000_101011101100;
            10'd0452: dout <= 36'b110100000110_000000011010_101011100001;
            10'd0453: dout <= 36'b110100001111_000000011100_101011010101;
            10'd0454: dout <= 36'b110100011001_000000011110_101011001001;
            10'd0455: dout <= 36'b110100100011_000000100000_101010111101;
            10'd0456: dout <= 36'b110100101100_000000100010_101010110010;
            10'd0457: dout <= 36'b110100110110_000000100100_101010100110;
            10'd0458: dout <= 36'b110100111111_000000100111_101010011010;
            10'd0459: dout <= 36'b110101001001_000000101001_101010001110;
            10'd0460: dout <= 36'b110101010010_000000101100_101010000010;
            10'd0461: dout <= 36'b110101011100_000000101110_101001110110;
            10'd0462: dout <= 36'b110101100101_000000110001_101001101010;
            10'd0463: dout <= 36'b110101101110_000000110100_101001011110;
            10'd0464: dout <= 36'b110101110111_000000110110_101001010010;
            10'd0465: dout <= 36'b110110000000_000000111001_101001000110;
            10'd0466: dout <= 36'b110110001010_000000111100_101000111010;
            10'd0467: dout <= 36'b110110010011_000000111111_101000101110;
            10'd0468: dout <= 36'b110110011100_000001000010_101000100010;
            10'd0469: dout <= 36'b110110100100_000001000110_101000010110;
            10'd0470: dout <= 36'b110110101101_000001001001_101000001010;
            10'd0471: dout <= 36'b110110110110_000001001100_100111111110;
            10'd0472: dout <= 36'b110110111111_000001010000_100111110001;
            10'd0473: dout <= 36'b110111001000_000001010011_100111100101;
            10'd0474: dout <= 36'b110111010000_000001010111_100111011001;
            10'd0475: dout <= 36'b110111011001_000001011010_100111001101;
            10'd0476: dout <= 36'b110111100001_000001011110_100111000001;
            10'd0477: dout <= 36'b110111101010_000001100010_100110110100;
            10'd0478: dout <= 36'b110111110010_000001100110_100110101000;
            10'd0479: dout <= 36'b110111111011_000001101010_100110011100;
            10'd0480: dout <= 36'b111000000011_000001101110_100110001111;
            10'd0481: dout <= 36'b111000001011_000001110010_100110000011;
            10'd0482: dout <= 36'b111000010011_000001110110_100101110111;
            10'd0483: dout <= 36'b111000011100_000001111010_100101101010;
            10'd0484: dout <= 36'b111000100100_000001111110_100101011110;
            10'd0485: dout <= 36'b111000101100_000010000011_100101010010;
            10'd0486: dout <= 36'b111000110100_000010000111_100101000101;
            10'd0487: dout <= 36'b111000111100_000010001100_100100111001;
            10'd0488: dout <= 36'b111001000011_000010010000_100100101100;
            10'd0489: dout <= 36'b111001001011_000010010101_100100100000;
            10'd0490: dout <= 36'b111001010011_000010011010_100100010011;
            10'd0491: dout <= 36'b111001011011_000010011110_100100000111;
            10'd0492: dout <= 36'b111001100010_000010100011_100011111011;
            10'd0493: dout <= 36'b111001101010_000010101000_100011101110;
            10'd0494: dout <= 36'b111001110001_000010101101_100011100010;
            10'd0495: dout <= 36'b111001111001_000010110010_100011010101;
            10'd0496: dout <= 36'b111010000000_000010110111_100011001001;
            10'd0497: dout <= 36'b111010000111_000010111101_100010111100;
            10'd0498: dout <= 36'b111010001110_000011000010_100010110000;
            10'd0499: dout <= 36'b111010010110_000011000111_100010100011;
            10'd0500: dout <= 36'b111010011101_000011001101_100010010111;
            10'd0501: dout <= 36'b111010100100_000011010010_100010001010;
            10'd0502: dout <= 36'b111010101011_000011011000_100001111110;
            10'd0503: dout <= 36'b111010110010_000011011101_100001110001;
            10'd0504: dout <= 36'b111010111000_000011100011_100001100100;
            10'd0505: dout <= 36'b111010111111_000011101001_100001011000;
            10'd0506: dout <= 36'b111011000110_000011101111_100001001011;
            10'd0507: dout <= 36'b111011001101_000011110101_100000111111;
            10'd0508: dout <= 36'b111011010011_000011111011_100000110010;
            10'd0509: dout <= 36'b111011011010_000100000001_100000100110;
            10'd0510: dout <= 36'b111011100000_000100000111_100000011001;
            10'd0511: dout <= 36'b111011100110_000100001101_100000001101;
            10'd0512: dout <= 36'b111011101101_000100010011_100000000000;
            10'd0513: dout <= 36'b111011110011_000100011010_011111110011;
            10'd0514: dout <= 36'b111011111001_000100100000_011111100111;
            10'd0515: dout <= 36'b111011111111_000100100110_011111011010;
            10'd0516: dout <= 36'b111100000101_000100101101_011111001110;
            10'd0517: dout <= 36'b111100001011_000100110011_011111000001;
            10'd0518: dout <= 36'b111100010001_000100111010_011110110101;
            10'd0519: dout <= 36'b111100010111_000101000001_011110101000;
            10'd0520: dout <= 36'b111100011101_000101001000_011110011100;
            10'd0521: dout <= 36'b111100100011_000101001110_011110001111;
            10'd0522: dout <= 36'b111100101000_000101010101_011110000010;
            10'd0523: dout <= 36'b111100101110_000101011100_011101110110;
            10'd0524: dout <= 36'b111100110011_000101100011_011101101001;
            10'd0525: dout <= 36'b111100111001_000101101010_011101011101;
            10'd0526: dout <= 36'b111100111110_000101110010_011101010000;
            10'd0527: dout <= 36'b111101000011_000101111001_011101000100;
            10'd0528: dout <= 36'b111101001001_000110000000_011100110111;
            10'd0529: dout <= 36'b111101001110_000110000111_011100101011;
            10'd0530: dout <= 36'b111101010011_000110001111_011100011110;
            10'd0531: dout <= 36'b111101011000_000110010110_011100010010;
            10'd0532: dout <= 36'b111101011101_000110011110_011100000101;
            10'd0533: dout <= 36'b111101100010_000110100101_011011111001;
            10'd0534: dout <= 36'b111101100110_000110101101_011011101101;
            10'd0535: dout <= 36'b111101101011_000110110101_011011100000;
            10'd0536: dout <= 36'b111101110000_000110111101_011011010100;
            10'd0537: dout <= 36'b111101110100_000111000100_011011000111;
            10'd0538: dout <= 36'b111101111001_000111001100_011010111011;
            10'd0539: dout <= 36'b111101111101_000111010100_011010101110;
            10'd0540: dout <= 36'b111110000010_000111011100_011010100010;
            10'd0541: dout <= 36'b111110000110_000111100100_011010010110;
            10'd0542: dout <= 36'b111110001010_000111101101_011010001001;
            10'd0543: dout <= 36'b111110001110_000111110101_011001111101;
            10'd0544: dout <= 36'b111110010010_000111111101_011001110001;
            10'd0545: dout <= 36'b111110010110_001000000101_011001100100;
            10'd0546: dout <= 36'b111110011010_001000001110_011001011000;
            10'd0547: dout <= 36'b111110011110_001000010110_011001001100;
            10'd0548: dout <= 36'b111110100010_001000011111_011000111111;
            10'd0549: dout <= 36'b111110100110_001000100111_011000110011;
            10'd0550: dout <= 36'b111110101001_001000110000_011000100111;
            10'd0551: dout <= 36'b111110101101_001000111000_011000011011;
            10'd0552: dout <= 36'b111110110000_001001000001_011000001111;
            10'd0553: dout <= 36'b111110110100_001001001010_011000000010;
            10'd0554: dout <= 36'b111110110111_001001010011_010111110110;
            10'd0555: dout <= 36'b111110111010_001001011100_010111101010;
            10'd0556: dout <= 36'b111110111110_001001100100_010111011110;
            10'd0557: dout <= 36'b111111000001_001001101101_010111010010;
            10'd0558: dout <= 36'b111111000100_001001110110_010111000110;
            10'd0559: dout <= 36'b111111000111_001010000000_010110111010;
            10'd0560: dout <= 36'b111111001010_001010001001_010110101110;
            10'd0561: dout <= 36'b111111001100_001010010010_010110100010;
            10'd0562: dout <= 36'b111111001111_001010011011_010110010110;
            10'd0563: dout <= 36'b111111010010_001010100100_010110001010;
            10'd0564: dout <= 36'b111111010100_001010101110_010101111110;
            10'd0565: dout <= 36'b111111010111_001010110111_010101110010;
            10'd0566: dout <= 36'b111111011001_001011000001_010101100110;
            10'd0567: dout <= 36'b111111011100_001011001010_010101011010;
            10'd0568: dout <= 36'b111111011110_001011010100_010101001110;
            10'd0569: dout <= 36'b111111100000_001011011101_010101000011;
            10'd0570: dout <= 36'b111111100010_001011100111_010100110111;
            10'd0571: dout <= 36'b111111100100_001011110001_010100101011;
            10'd0572: dout <= 36'b111111100110_001011111010_010100011111;
            10'd0573: dout <= 36'b111111101000_001100000100_010100010100;
            10'd0574: dout <= 36'b111111101010_001100001110_010100001000;
            10'd0575: dout <= 36'b111111101100_001100011000_010011111100;
            10'd0576: dout <= 36'b111111101101_001100100010_010011110001;
            10'd0577: dout <= 36'b111111101111_001100101100_010011100101;
            10'd0578: dout <= 36'b111111110001_001100110110_010011011001;
            10'd0579: dout <= 36'b111111110010_001101000000_010011001110;
            10'd0580: dout <= 36'b111111110011_001101001010_010011000010;
            10'd0581: dout <= 36'b111111110101_001101010100_010010110111;
            10'd0582: dout <= 36'b111111110110_001101011110_010010101100;
            10'd0583: dout <= 36'b111111110111_001101101001_010010100000;
            10'd0584: dout <= 36'b111111111000_001101110011_010010010101;
            10'd0585: dout <= 36'b111111111001_001101111101_010010001001;
            10'd0586: dout <= 36'b111111111010_001110001000_010001111110;
            10'd0587: dout <= 36'b111111111011_001110010010_010001110011;
            10'd0588: dout <= 36'b111111111100_001110011101_010001101000;
            10'd0589: dout <= 36'b111111111100_001110100111_010001011100;
            10'd0590: dout <= 36'b111111111101_001110110010_010001010001;
            10'd0591: dout <= 36'b111111111101_001110111100_010001000110;
            10'd0592: dout <= 36'b111111111110_001111000111_010000111011;
            10'd0593: dout <= 36'b111111111110_001111010010_010000110000;
            10'd0594: dout <= 36'b111111111111_001111011100_010000100101;
            10'd0595: dout <= 36'b111111111111_001111100111_010000011010;
            10'd0596: dout <= 36'b111111111111_001111110010_010000001111;
            10'd0597: dout <= 36'b111111111111_001111111101_010000000100;
            10'd0598: dout <= 36'b111111111111_010000001000_001111111001;
            10'd0599: dout <= 36'b111111111111_010000010011_001111101110;
            10'd0600: dout <= 36'b111111111111_010000011110_001111100100;
            10'd0601: dout <= 36'b111111111110_010000101001_001111011001;
            10'd0602: dout <= 36'b111111111110_010000110100_001111001110;
            10'd0603: dout <= 36'b111111111110_010000111111_001111000011;
            10'd0604: dout <= 36'b111111111101_010001001010_001110111001;
            10'd0605: dout <= 36'b111111111101_010001010101_001110101110;
            10'd0606: dout <= 36'b111111111100_010001100000_001110100100;
            10'd0607: dout <= 36'b111111111011_010001101011_001110011001;
            10'd0608: dout <= 36'b111111111011_010001110111_001110001111;
            10'd0609: dout <= 36'b111111111010_010010000010_001110000100;
            10'd0610: dout <= 36'b111111111001_010010001101_001101111010;
            10'd0611: dout <= 36'b111111111000_010010011001_001101110000;
            10'd0612: dout <= 36'b111111110111_010010100100_001101100101;
            10'd0613: dout <= 36'b111111110110_010010101111_001101011011;
            10'd0614: dout <= 36'b111111110100_010010111011_001101010001;
            10'd0615: dout <= 36'b111111110011_010011000110_001101000111;
            10'd0616: dout <= 36'b111111110010_010011010010_001100111101;
            10'd0617: dout <= 36'b111111110000_010011011101_001100110011;
            10'd0618: dout <= 36'b111111101111_010011101001_001100101001;
            10'd0619: dout <= 36'b111111101101_010011110101_001100011111;
            10'd0620: dout <= 36'b111111101011_010100000000_001100010101;
            10'd0621: dout <= 36'b111111101001_010100001100_001100001011;
            10'd0622: dout <= 36'b111111101000_010100010111_001100000001;
            10'd0623: dout <= 36'b111111100110_010100100011_001011110111;
            10'd0624: dout <= 36'b111111100100_010100101111_001011101101;
            10'd0625: dout <= 36'b111111100010_010100111011_001011100100;
            10'd0626: dout <= 36'b111111011111_010101000111_001011011010;
            10'd0627: dout <= 36'b111111011101_010101010010_001011010000;
            10'd0628: dout <= 36'b111111011011_010101011110_001011000111;
            10'd0629: dout <= 36'b111111011000_010101101010_001010111101;
            10'd0630: dout <= 36'b111111010110_010101110110_001010110100;
            10'd0631: dout <= 36'b111111010011_010110000010_001010101011;
            10'd0632: dout <= 36'b111111010001_010110001110_001010100001;
            10'd0633: dout <= 36'b111111001110_010110011010_001010011000;
            10'd0634: dout <= 36'b111111001011_010110100110_001010001111;
            10'd0635: dout <= 36'b111111001001_010110110010_001010000110;
            10'd0636: dout <= 36'b111111000110_010110111110_001001111101;
            10'd0637: dout <= 36'b111111000011_010111001010_001001110011;
            10'd0638: dout <= 36'b111111000000_010111010110_001001101010;
            10'd0639: dout <= 36'b111110111100_010111100010_001001100001;
            10'd0640: dout <= 36'b111110111001_010111101110_001001011001;
            10'd0641: dout <= 36'b111110110110_010111111010_001001010000;
            10'd0642: dout <= 36'b111110110011_011000000111_001001000111;
            10'd0643: dout <= 36'b111110101111_011000010011_001000111110;
            10'd0644: dout <= 36'b111110101100_011000011111_001000110101;
            10'd0645: dout <= 36'b111110101000_011000101011_001000101101;
            10'd0646: dout <= 36'b111110100100_011000110111_001000100100;
            10'd0647: dout <= 36'b111110100001_011001000100_001000011100;
            10'd0648: dout <= 36'b111110011101_011001010000_001000010011;
            10'd0649: dout <= 36'b111110011001_011001011100_001000001011;
            10'd0650: dout <= 36'b111110010101_011001101000_001000000011;
            10'd0651: dout <= 36'b111110010001_011001110101_000111111010;
            10'd0652: dout <= 36'b111110001101_011010000001_000111110010;
            10'd0653: dout <= 36'b111110001001_011010001101_000111101010;
            10'd0654: dout <= 36'b111110000101_011010011010_000111100010;
            10'd0655: dout <= 36'b111110000000_011010100110_000111011010;
            10'd0656: dout <= 36'b111101111100_011010110011_000111010010;
            10'd0657: dout <= 36'b111101110111_011010111111_000111001010;
            10'd0658: dout <= 36'b111101110011_011011001011_000111000010;
            10'd0659: dout <= 36'b111101101110_011011011000_000110111010;
            10'd0660: dout <= 36'b111101101010_011011100100_000110110010;
            10'd0661: dout <= 36'b111101100101_011011110001_000110101011;
            10'd0662: dout <= 36'b111101100000_011011111101_000110100011;
            10'd0663: dout <= 36'b111101011011_011100001010_000110011011;
            10'd0664: dout <= 36'b111101010110_011100010110_000110010100;
            10'd0665: dout <= 36'b111101010001_011100100011_000110001100;
            10'd0666: dout <= 36'b111101001100_011100101111_000110000101;
            10'd0667: dout <= 36'b111101000111_011100111100_000101111110;
            10'd0668: dout <= 36'b111101000010_011101001000_000101110110;
            10'd0669: dout <= 36'b111100111100_011101010101_000101101111;
            10'd0670: dout <= 36'b111100110111_011101100001_000101101000;
            10'd0671: dout <= 36'b111100110001_011101101110_000101100001;
            10'd0672: dout <= 36'b111100101100_011101111010_000101011010;
            10'd0673: dout <= 36'b111100100110_011110000111_000101010011;
            10'd0674: dout <= 36'b111100100001_011110010011_000101001100;
            10'd0675: dout <= 36'b111100011011_011110100000_000101000101;
            10'd0676: dout <= 36'b111100010101_011110101100_000100111111;
            10'd0677: dout <= 36'b111100001111_011110111001_000100111000;
            10'd0678: dout <= 36'b111100001001_011111000101_000100110001;
            10'd0679: dout <= 36'b111100000011_011111010010_000100101011;
            10'd0680: dout <= 36'b111011111101_011111011111_000100100100;
            10'd0681: dout <= 36'b111011110111_011111101011_000100011110;
            10'd0682: dout <= 36'b111011110001_011111111000_000100010111;
            10'd0683: dout <= 36'b111011101011_100000000100_000100010001;
            10'd0684: dout <= 36'b111011100100_100000010001_000100001011;
            10'd0685: dout <= 36'b111011011110_100000011101_000100000101;
            10'd0686: dout <= 36'b111011010111_100000101010_000011111111;
            10'd0687: dout <= 36'b111011010001_100000110110_000011111001;
            10'd0688: dout <= 36'b111011001010_100001000011_000011110011;
            10'd0689: dout <= 36'b111011000100_100001010000_000011101101;
            10'd0690: dout <= 36'b111010111101_100001011100_000011100111;
            10'd0691: dout <= 36'b111010110110_100001101001_000011100001;
            10'd0692: dout <= 36'b111010101111_100001110101_000011011100;
            10'd0693: dout <= 36'b111010101000_100010000010_000011010110;
            10'd0694: dout <= 36'b111010100001_100010001110_000011010000;
            10'd0695: dout <= 36'b111010011010_100010011011_000011001011;
            10'd0696: dout <= 36'b111010010011_100010100111_000011000110;
            10'd0697: dout <= 36'b111010001100_100010110100_000011000000;
            10'd0698: dout <= 36'b111010000101_100011000000_000010111011;
            10'd0699: dout <= 36'b111001111101_100011001101_000010110110;
            10'd0700: dout <= 36'b111001110110_100011011001_000010110001;
            10'd0701: dout <= 36'b111001101111_100011100110_000010101100;
            10'd0702: dout <= 36'b111001100111_100011110010_000010100111;
            10'd0703: dout <= 36'b111001100000_100011111111_000010100010;
            10'd0704: dout <= 36'b111001011000_100100001011_000010011101;
            10'd0705: dout <= 36'b111001010000_100100011000_000010011000;
            10'd0706: dout <= 36'b111001001001_100100100100_000010010011;
            10'd0707: dout <= 36'b111001000001_100100110000_000010001111;
            10'd0708: dout <= 36'b111000111001_100100111101_000010001010;
            10'd0709: dout <= 36'b111000110001_100101001001_000010000110;
            10'd0710: dout <= 36'b111000101001_100101010110_000010000001;
            10'd0711: dout <= 36'b111000100001_100101100010_000001111101;
            10'd0712: dout <= 36'b111000011001_100101101110_000001111001;
            10'd0713: dout <= 36'b111000010001_100101111011_000001110100;
            10'd0714: dout <= 36'b111000001001_100110000111_000001110000;
            10'd0715: dout <= 36'b111000000000_100110010011_000001101100;
            10'd0716: dout <= 36'b110111111000_100110100000_000001101000;
            10'd0717: dout <= 36'b110111110000_100110101100_000001100100;
            10'd0718: dout <= 36'b110111100111_100110111000_000001100001;
            10'd0719: dout <= 36'b110111011111_100111000101_000001011101;
            10'd0720: dout <= 36'b110111010110_100111010001_000001011001;
            10'd0721: dout <= 36'b110111001101_100111011101_000001010110;
            10'd0722: dout <= 36'b110111000101_100111101001_000001010010;
            10'd0723: dout <= 36'b110110111100_100111110101_000001001111;
            10'd0724: dout <= 36'b110110110011_101000000010_000001001011;
            10'd0725: dout <= 36'b110110101010_101000001110_000001001000;
            10'd0726: dout <= 36'b110110100010_101000011010_000001000101;
            10'd0727: dout <= 36'b110110011001_101000100110_000001000001;
            10'd0728: dout <= 36'b110110010000_101000110010_000000111110;
            10'd0729: dout <= 36'b110110000111_101000111110_000000111011;
            10'd0730: dout <= 36'b110101111101_101001001010_000000111000;
            10'd0731: dout <= 36'b110101110100_101001010110_000000110110;
            10'd0732: dout <= 36'b110101101011_101001100010_000000110011;
            10'd0733: dout <= 36'b110101100010_101001101110_000000110000;
            10'd0734: dout <= 36'b110101011000_101001111010_000000101101;
            10'd0735: dout <= 36'b110101001111_101010000110_000000101011;
            10'd0736: dout <= 36'b110101000110_101010010010_000000101000;
            10'd0737: dout <= 36'b110100111100_101010011110_000000100110;
            10'd0738: dout <= 36'b110100110011_101010101010_000000100100;
            10'd0739: dout <= 36'b110100101001_101010110110_000000100001;
            10'd0740: dout <= 36'b110100100000_101011000001_000000011111;
            10'd0741: dout <= 36'b110100010110_101011001101_000000011101;
            10'd0742: dout <= 36'b110100001100_101011011001_000000011011;
            10'd0743: dout <= 36'b110100000010_101011100101_000000011001;
            10'd0744: dout <= 36'b110011111001_101011110000_000000010111;
            10'd0745: dout <= 36'b110011101111_101011111100_000000010101;
            10'd0746: dout <= 36'b110011100101_101100001000_000000010100;
            10'd0747: dout <= 36'b110011011011_101100010011_000000010010;
            10'd0748: dout <= 36'b110011010001_101100011111_000000010000;
            10'd0749: dout <= 36'b110011000111_101100101010_000000001111;
            10'd0750: dout <= 36'b110010111101_101100110110_000000001101;
            10'd0751: dout <= 36'b110010110011_101101000001_000000001100;
            10'd0752: dout <= 36'b110010101000_101101001101_000000001011;
            10'd0753: dout <= 36'b110010011110_101101011000_000000001010;
            10'd0754: dout <= 36'b110010010100_101101100100_000000001001;
            10'd0755: dout <= 36'b110010001010_101101101111_000000001000;
            10'd0756: dout <= 36'b110001111111_101101111010_000000000111;
            10'd0757: dout <= 36'b110001110101_101110000110_000000000110;
            10'd0758: dout <= 36'b110001101010_101110010001_000000000101;
            10'd0759: dout <= 36'b110001100000_101110011100_000000000100;
            10'd0760: dout <= 36'b110001010101_101110100111_000000000011;
            10'd0761: dout <= 36'b110001001011_101110110010_000000000011;
            10'd0762: dout <= 36'b110001000000_101110111110_000000000010;
            10'd0763: dout <= 36'b110000110101_101111001001_000000000010;
            10'd0764: dout <= 36'b110000101011_101111010100_000000000010;
            10'd0765: dout <= 36'b110000100000_101111011111_000000000001;
            10'd0766: dout <= 36'b110000010101_101111101010_000000000001;
            10'd0767: dout <= 36'b110000001010_101111110101_000000000001;
            10'd0768: dout <= 36'b101111111111_101111111111_000000000001;
            10'd0769: dout <= 36'b101111110101_110000001010_000000000001;
            10'd0770: dout <= 36'b101111101010_110000010101_000000000001;
            10'd0771: dout <= 36'b101111011111_110000100000_000000000001;
            10'd0772: dout <= 36'b101111010100_110000101011_000000000010;
            10'd0773: dout <= 36'b101111001001_110000110101_000000000010;
            10'd0774: dout <= 36'b101110111110_110001000000_000000000010;
            10'd0775: dout <= 36'b101110110010_110001001011_000000000011;
            10'd0776: dout <= 36'b101110100111_110001010101_000000000011;
            10'd0777: dout <= 36'b101110011100_110001100000_000000000100;
            10'd0778: dout <= 36'b101110010001_110001101010_000000000101;
            10'd0779: dout <= 36'b101110000110_110001110101_000000000110;
            10'd0780: dout <= 36'b101101111010_110001111111_000000000111;
            10'd0781: dout <= 36'b101101101111_110010001010_000000001000;
            10'd0782: dout <= 36'b101101100100_110010010100_000000001001;
            10'd0783: dout <= 36'b101101011000_110010011110_000000001010;
            10'd0784: dout <= 36'b101101001101_110010101000_000000001011;
            10'd0785: dout <= 36'b101101000001_110010110011_000000001100;
            10'd0786: dout <= 36'b101100110110_110010111101_000000001101;
            10'd0787: dout <= 36'b101100101010_110011000111_000000001111;
            10'd0788: dout <= 36'b101100011111_110011010001_000000010000;
            10'd0789: dout <= 36'b101100010011_110011011011_000000010010;
            10'd0790: dout <= 36'b101100001000_110011100101_000000010100;
            10'd0791: dout <= 36'b101011111100_110011101111_000000010101;
            10'd0792: dout <= 36'b101011110000_110011111001_000000010111;
            10'd0793: dout <= 36'b101011100101_110100000010_000000011001;
            10'd0794: dout <= 36'b101011011001_110100001100_000000011011;
            10'd0795: dout <= 36'b101011001101_110100010110_000000011101;
            10'd0796: dout <= 36'b101011000001_110100100000_000000011111;
            10'd0797: dout <= 36'b101010110110_110100101001_000000100001;
            10'd0798: dout <= 36'b101010101010_110100110011_000000100100;
            10'd0799: dout <= 36'b101010011110_110100111100_000000100110;
            10'd0800: dout <= 36'b101010010010_110101000110_000000101000;
            10'd0801: dout <= 36'b101010000110_110101001111_000000101011;
            10'd0802: dout <= 36'b101001111010_110101011000_000000101101;
            10'd0803: dout <= 36'b101001101110_110101100010_000000110000;
            10'd0804: dout <= 36'b101001100010_110101101011_000000110011;
            10'd0805: dout <= 36'b101001010110_110101110100_000000110110;
            10'd0806: dout <= 36'b101001001010_110101111101_000000111000;
            10'd0807: dout <= 36'b101000111110_110110000111_000000111011;
            10'd0808: dout <= 36'b101000110010_110110010000_000000111110;
            10'd0809: dout <= 36'b101000100110_110110011001_000001000001;
            10'd0810: dout <= 36'b101000011010_110110100010_000001000101;
            10'd0811: dout <= 36'b101000001110_110110101010_000001001000;
            10'd0812: dout <= 36'b101000000010_110110110011_000001001011;
            10'd0813: dout <= 36'b100111110101_110110111100_000001001111;
            10'd0814: dout <= 36'b100111101001_110111000101_000001010010;
            10'd0815: dout <= 36'b100111011101_110111001101_000001010110;
            10'd0816: dout <= 36'b100111010001_110111010110_000001011001;
            10'd0817: dout <= 36'b100111000101_110111011111_000001011101;
            10'd0818: dout <= 36'b100110111000_110111100111_000001100001;
            10'd0819: dout <= 36'b100110101100_110111110000_000001100100;
            10'd0820: dout <= 36'b100110100000_110111111000_000001101000;
            10'd0821: dout <= 36'b100110010011_111000000000_000001101100;
            10'd0822: dout <= 36'b100110000111_111000001001_000001110000;
            10'd0823: dout <= 36'b100101111011_111000010001_000001110100;
            10'd0824: dout <= 36'b100101101110_111000011001_000001111001;
            10'd0825: dout <= 36'b100101100010_111000100001_000001111101;
            10'd0826: dout <= 36'b100101010110_111000101001_000010000001;
            10'd0827: dout <= 36'b100101001001_111000110001_000010000110;
            10'd0828: dout <= 36'b100100111101_111000111001_000010001010;
            10'd0829: dout <= 36'b100100110000_111001000001_000010001111;
            10'd0830: dout <= 36'b100100100100_111001001001_000010010011;
            10'd0831: dout <= 36'b100100011000_111001010000_000010011000;
            10'd0832: dout <= 36'b100100001011_111001011000_000010011101;
            10'd0833: dout <= 36'b100011111111_111001100000_000010100010;
            10'd0834: dout <= 36'b100011110010_111001100111_000010100111;
            10'd0835: dout <= 36'b100011100110_111001101111_000010101100;
            10'd0836: dout <= 36'b100011011001_111001110110_000010110001;
            10'd0837: dout <= 36'b100011001101_111001111101_000010110110;
            10'd0838: dout <= 36'b100011000000_111010000101_000010111011;
            10'd0839: dout <= 36'b100010110100_111010001100_000011000000;
            10'd0840: dout <= 36'b100010100111_111010010011_000011000110;
            10'd0841: dout <= 36'b100010011011_111010011010_000011001011;
            10'd0842: dout <= 36'b100010001110_111010100001_000011010000;
            10'd0843: dout <= 36'b100010000010_111010101000_000011010110;
            10'd0844: dout <= 36'b100001110101_111010101111_000011011100;
            10'd0845: dout <= 36'b100001101001_111010110110_000011100001;
            10'd0846: dout <= 36'b100001011100_111010111101_000011100111;
            10'd0847: dout <= 36'b100001010000_111011000100_000011101101;
            10'd0848: dout <= 36'b100001000011_111011001010_000011110011;
            10'd0849: dout <= 36'b100000110110_111011010001_000011111001;
            10'd0850: dout <= 36'b100000101010_111011010111_000011111111;
            10'd0851: dout <= 36'b100000011101_111011011110_000100000101;
            10'd0852: dout <= 36'b100000010001_111011100100_000100001011;
            10'd0853: dout <= 36'b100000000100_111011101011_000100010001;
            10'd0854: dout <= 36'b011111111000_111011110001_000100010111;
            10'd0855: dout <= 36'b011111101011_111011110111_000100011110;
            10'd0856: dout <= 36'b011111011111_111011111101_000100100100;
            10'd0857: dout <= 36'b011111010010_111100000011_000100101011;
            10'd0858: dout <= 36'b011111000101_111100001001_000100110001;
            10'd0859: dout <= 36'b011110111001_111100001111_000100111000;
            10'd0860: dout <= 36'b011110101100_111100010101_000100111111;
            10'd0861: dout <= 36'b011110100000_111100011011_000101000101;
            10'd0862: dout <= 36'b011110010011_111100100001_000101001100;
            10'd0863: dout <= 36'b011110000111_111100100110_000101010011;
            10'd0864: dout <= 36'b011101111010_111100101100_000101011010;
            10'd0865: dout <= 36'b011101101110_111100110001_000101100001;
            10'd0866: dout <= 36'b011101100001_111100110111_000101101000;
            10'd0867: dout <= 36'b011101010101_111100111100_000101101111;
            10'd0868: dout <= 36'b011101001000_111101000010_000101110110;
            10'd0869: dout <= 36'b011100111100_111101000111_000101111110;
            10'd0870: dout <= 36'b011100101111_111101001100_000110000101;
            10'd0871: dout <= 36'b011100100011_111101010001_000110001100;
            10'd0872: dout <= 36'b011100010110_111101010110_000110010100;
            10'd0873: dout <= 36'b011100001010_111101011011_000110011011;
            10'd0874: dout <= 36'b011011111101_111101100000_000110100011;
            10'd0875: dout <= 36'b011011110001_111101100101_000110101011;
            10'd0876: dout <= 36'b011011100100_111101101010_000110110010;
            10'd0877: dout <= 36'b011011011000_111101101110_000110111010;
            10'd0878: dout <= 36'b011011001011_111101110011_000111000010;
            10'd0879: dout <= 36'b011010111111_111101110111_000111001010;
            10'd0880: dout <= 36'b011010110011_111101111100_000111010010;
            10'd0881: dout <= 36'b011010100110_111110000000_000111011010;
            10'd0882: dout <= 36'b011010011010_111110000101_000111100010;
            10'd0883: dout <= 36'b011010001101_111110001001_000111101010;
            10'd0884: dout <= 36'b011010000001_111110001101_000111110010;
            10'd0885: dout <= 36'b011001110101_111110010001_000111111010;
            10'd0886: dout <= 36'b011001101000_111110010101_001000000011;
            10'd0887: dout <= 36'b011001011100_111110011001_001000001011;
            10'd0888: dout <= 36'b011001010000_111110011101_001000010011;
            10'd0889: dout <= 36'b011001000100_111110100001_001000011100;
            10'd0890: dout <= 36'b011000110111_111110100100_001000100100;
            10'd0891: dout <= 36'b011000101011_111110101000_001000101101;
            10'd0892: dout <= 36'b011000011111_111110101100_001000110101;
            10'd0893: dout <= 36'b011000010011_111110101111_001000111110;
            10'd0894: dout <= 36'b011000000111_111110110011_001001000111;
            10'd0895: dout <= 36'b010111111010_111110110110_001001010000;
            10'd0896: dout <= 36'b010111101110_111110111001_001001011001;
            10'd0897: dout <= 36'b010111100010_111110111100_001001100001;
            10'd0898: dout <= 36'b010111010110_111111000000_001001101010;
            10'd0899: dout <= 36'b010111001010_111111000011_001001110011;
            10'd0900: dout <= 36'b010110111110_111111000110_001001111101;
            10'd0901: dout <= 36'b010110110010_111111001001_001010000110;
            10'd0902: dout <= 36'b010110100110_111111001011_001010001111;
            10'd0903: dout <= 36'b010110011010_111111001110_001010011000;
            10'd0904: dout <= 36'b010110001110_111111010001_001010100001;
            10'd0905: dout <= 36'b010110000010_111111010011_001010101011;
            10'd0906: dout <= 36'b010101110110_111111010110_001010110100;
            10'd0907: dout <= 36'b010101101010_111111011000_001010111101;
            10'd0908: dout <= 36'b010101011110_111111011011_001011000111;
            10'd0909: dout <= 36'b010101010010_111111011101_001011010000;
            10'd0910: dout <= 36'b010101000111_111111011111_001011011010;
            10'd0911: dout <= 36'b010100111011_111111100010_001011100100;
            10'd0912: dout <= 36'b010100101111_111111100100_001011101101;
            10'd0913: dout <= 36'b010100100011_111111100110_001011110111;
            10'd0914: dout <= 36'b010100010111_111111101000_001100000001;
            10'd0915: dout <= 36'b010100001100_111111101001_001100001011;
            10'd0916: dout <= 36'b010100000000_111111101011_001100010101;
            10'd0917: dout <= 36'b010011110101_111111101101_001100011111;
            10'd0918: dout <= 36'b010011101001_111111101111_001100101001;
            10'd0919: dout <= 36'b010011011101_111111110000_001100110011;
            10'd0920: dout <= 36'b010011010010_111111110010_001100111101;
            10'd0921: dout <= 36'b010011000110_111111110011_001101000111;
            10'd0922: dout <= 36'b010010111011_111111110100_001101010001;
            10'd0923: dout <= 36'b010010101111_111111110110_001101011011;
            10'd0924: dout <= 36'b010010100100_111111110111_001101100101;
            10'd0925: dout <= 36'b010010011001_111111111000_001101110000;
            10'd0926: dout <= 36'b010010001101_111111111001_001101111010;
            10'd0927: dout <= 36'b010010000010_111111111010_001110000100;
            10'd0928: dout <= 36'b010001110111_111111111011_001110001111;
            10'd0929: dout <= 36'b010001101011_111111111011_001110011001;
            10'd0930: dout <= 36'b010001100000_111111111100_001110100100;
            10'd0931: dout <= 36'b010001010101_111111111101_001110101110;
            10'd0932: dout <= 36'b010001001010_111111111101_001110111001;
            10'd0933: dout <= 36'b010000111111_111111111110_001111000011;
            10'd0934: dout <= 36'b010000110100_111111111110_001111001110;
            10'd0935: dout <= 36'b010000101001_111111111110_001111011001;
            10'd0936: dout <= 36'b010000011110_111111111111_001111100100;
            10'd0937: dout <= 36'b010000010011_111111111111_001111101110;
            10'd0938: dout <= 36'b010000001000_111111111111_001111111001;
            10'd0939: dout <= 36'b001111111101_111111111111_010000000100;
            10'd0940: dout <= 36'b001111110010_111111111111_010000001111;
            10'd0941: dout <= 36'b001111100111_111111111111_010000011010;
            10'd0942: dout <= 36'b001111011100_111111111111_010000100101;
            10'd0943: dout <= 36'b001111010010_111111111110_010000110000;
            10'd0944: dout <= 36'b001111000111_111111111110_010000111011;
            10'd0945: dout <= 36'b001110111100_111111111101_010001000110;
            10'd0946: dout <= 36'b001110110010_111111111101_010001010001;
            10'd0947: dout <= 36'b001110100111_111111111100_010001011100;
            10'd0948: dout <= 36'b001110011101_111111111100_010001101000;
            10'd0949: dout <= 36'b001110010010_111111111011_010001110011;
            10'd0950: dout <= 36'b001110001000_111111111010_010001111110;
            10'd0951: dout <= 36'b001101111101_111111111001_010010001001;
            10'd0952: dout <= 36'b001101110011_111111111000_010010010101;
            10'd0953: dout <= 36'b001101101001_111111110111_010010100000;
            10'd0954: dout <= 36'b001101011110_111111110110_010010101100;
            10'd0955: dout <= 36'b001101010100_111111110101_010010110111;
            10'd0956: dout <= 36'b001101001010_111111110011_010011000010;
            10'd0957: dout <= 36'b001101000000_111111110010_010011001110;
            10'd0958: dout <= 36'b001100110110_111111110001_010011011001;
            10'd0959: dout <= 36'b001100101100_111111101111_010011100101;
            10'd0960: dout <= 36'b001100100010_111111101101_010011110001;
            10'd0961: dout <= 36'b001100011000_111111101100_010011111100;
            10'd0962: dout <= 36'b001100001110_111111101010_010100001000;
            10'd0963: dout <= 36'b001100000100_111111101000_010100010100;
            10'd0964: dout <= 36'b001011111010_111111100110_010100011111;
            10'd0965: dout <= 36'b001011110001_111111100100_010100101011;
            10'd0966: dout <= 36'b001011100111_111111100010_010100110111;
            10'd0967: dout <= 36'b001011011101_111111100000_010101000011;
            10'd0968: dout <= 36'b001011010100_111111011110_010101001110;
            10'd0969: dout <= 36'b001011001010_111111011100_010101011010;
            10'd0970: dout <= 36'b001011000001_111111011001_010101100110;
            10'd0971: dout <= 36'b001010110111_111111010111_010101110010;
            10'd0972: dout <= 36'b001010101110_111111010100_010101111110;
            10'd0973: dout <= 36'b001010100100_111111010010_010110001010;
            10'd0974: dout <= 36'b001010011011_111111001111_010110010110;
            10'd0975: dout <= 36'b001010010010_111111001100_010110100010;
            10'd0976: dout <= 36'b001010001001_111111001010_010110101110;
            10'd0977: dout <= 36'b001010000000_111111000111_010110111010;
            10'd0978: dout <= 36'b001001110110_111111000100_010111000110;
            10'd0979: dout <= 36'b001001101101_111111000001_010111010010;
            10'd0980: dout <= 36'b001001100100_111110111110_010111011110;
            10'd0981: dout <= 36'b001001011100_111110111010_010111101010;
            10'd0982: dout <= 36'b001001010011_111110110111_010111110110;
            10'd0983: dout <= 36'b001001001010_111110110100_011000000010;
            10'd0984: dout <= 36'b001001000001_111110110000_011000001111;
            10'd0985: dout <= 36'b001000111000_111110101101_011000011011;
            10'd0986: dout <= 36'b001000110000_111110101001_011000100111;
            10'd0987: dout <= 36'b001000100111_111110100110_011000110011;
            10'd0988: dout <= 36'b001000011111_111110100010_011000111111;
            10'd0989: dout <= 36'b001000010110_111110011110_011001001100;
            10'd0990: dout <= 36'b001000001110_111110011010_011001011000;
            10'd0991: dout <= 36'b001000000101_111110010110_011001100100;
            10'd0992: dout <= 36'b000111111101_111110010010_011001110001;
            10'd0993: dout <= 36'b000111110101_111110001110_011001111101;
            10'd0994: dout <= 36'b000111101101_111110001010_011010001001;
            10'd0995: dout <= 36'b000111100100_111110000110_011010010110;
            10'd0996: dout <= 36'b000111011100_111110000010_011010100010;
            10'd0997: dout <= 36'b000111010100_111101111101_011010101110;
            10'd0998: dout <= 36'b000111001100_111101111001_011010111011;
            10'd0999: dout <= 36'b000111000100_111101110100_011011000111;
            10'd1000: dout <= 36'b000110111101_111101110000_011011010100;
            10'd1001: dout <= 36'b000110110101_111101101011_011011100000;
            10'd1002: dout <= 36'b000110101101_111101100110_011011101101;
            10'd1003: dout <= 36'b000110100101_111101100010_011011111001;
            10'd1004: dout <= 36'b000110011110_111101011101_011100000101;
            10'd1005: dout <= 36'b000110010110_111101011000_011100010010;
            10'd1006: dout <= 36'b000110001111_111101010011_011100011110;
            10'd1007: dout <= 36'b000110000111_111101001110_011100101011;
            10'd1008: dout <= 36'b000110000000_111101001001_011100110111;
            10'd1009: dout <= 36'b000101111001_111101000011_011101000100;
            10'd1010: dout <= 36'b000101110010_111100111110_011101010000;
            10'd1011: dout <= 36'b000101101010_111100111001_011101011101;
            10'd1012: dout <= 36'b000101100011_111100110011_011101101001;
            10'd1013: dout <= 36'b000101011100_111100101110_011101110110;
            10'd1014: dout <= 36'b000101010101_111100101000_011110000010;
            10'd1015: dout <= 36'b000101001110_111100100011_011110001111;
            10'd1016: dout <= 36'b000101001000_111100011101_011110011100;
            10'd1017: dout <= 36'b000101000001_111100010111_011110101000;
            10'd1018: dout <= 36'b000100111010_111100010001_011110110101;
            10'd1019: dout <= 36'b000100110011_111100001011_011111000001;
            10'd1020: dout <= 36'b000100101101_111100000101_011111001110;
            10'd1021: dout <= 36'b000100100110_111011111111_011111011010;
            10'd1022: dout <= 36'b000100100000_111011111001_011111100111;
            10'd1023: dout <= 36'b000100011010_111011110011_011111110011;
            endcase
        end
    end
    
    assign {out_z, out_y, out_x} = dout;
    
    
endmodule


`default_nettype wire


// end of file

