
`timescale 1 ns / 1 ps

module design_1
   (
    fan_en);
  output fan_en;
  wire fan_en;

  assign fan_en = 1'b0  ;

endmodule
