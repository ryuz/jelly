`timescale 1 ps / 1 ps

module kv260_axi_test
        (
            output   var logic   fan_en
        );
    
  design_1
    u_design_1
        (
            .fan_en (fan_en)
        );

endmodule

